`timescale 1ns / 1ps
module F_short_t12_next_Rom5(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[167:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 168'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h14: rd_q <= 168'b010000110100100101011011100100001101011111010000001110010000011001001101011101011001010001110100111010100101000111011101000101010111111101001011101010000001000111110001;
			5'h13: rd_q <= 168'b011111111001110101100110110010011101011101010101001001001010011000101001010101111011101110100010101011010110010001011010100001000000001101111001010000011011011000101100;
			5'h12: rd_q <= 168'b010010010110110011001111011111101010000010111001000100110011011001000010001111000101111110010011000000111100100011011101100101101001101011011101101011001110010000100111;
			5'h11: rd_q <= 168'b000010011100111010100110000101001111100001100110100101100010000000100000010101101001010010011111010000111001110000111001101010011000001101011000010100001100001100010000;
			5'h10: rd_q <= 168'b010001100110110110010001111100101001110001110111011000000001101000111001111001011000110011001110010100001000100001110011010000000110011000000010010011101001101100000010;
			5'h0f: rd_q <= 168'b100001000100001001011000110100100111001010010011100110101010100110101010100010101110101001110010000010000011111000101011011011111110011010010100000011010000000001100001;
			5'h0e: rd_q <= 168'b100111001001111010101010000101011111011010011000100100001100001100001001011111000101101101000010110101110000101110010111100111011010111100110110010100111001111011111110;
			5'h0d: rd_q <= 168'b011111001001111101110010011010110110101000001100001111000010100001010011011001111000011011110001000000001111001010010101011000111111111111111110110011001001011000110111;
			5'h0c: rd_q <= 168'b010011111001111100001010111111010110010100100011001001011000001100100111100000100001010100011100111011100101010011101100100110001011100110111100011001010110100010100011;
			5'h0b: rd_q <= 168'b111011110010000110010110110010100100011110010100110001000101101001001110010011110111101101100101100101010110011000110101000110111110101101100111010000100101110101101111;
			5'h0a: rd_q <= 168'b110111010010101000010000001010010001011011010010001100010101111010011101101101010010110110110000001110000000101000001011101000001111110000010101010101111010110101001010;
			5'h09: rd_q <= 168'b010100001001101111100100001101111111001101001010101101010101000100111111110000010111000011011000111110110101011000110101111101101111010000110010101001111001100110110100;
			5'h08: rd_q <= 168'b001011000001010110111001000000101001001001010101100010010110110110100000000011011111111000101111110100011011000011110111001111001100000001101011011110101010110000101001;
			5'h07: rd_q <= 168'b010010000111010000000110100100000111110000101011110111000111100100011100100110010001011001011101000001111101001010000101101000000000111000101100000100010110100110110001;
			5'h06: rd_q <= 168'b001011010100011000010111110100010010001000001101001001111110011000011101000000101011010111000010110111010010101011111111000101111011101010100011110010111010110001010101;
			5'h05: rd_q <= 168'b000101011101001000010100001101111011101110001001001111001110110000100001111100000010100110000110110111011101001101101111110101101111100010100010111101110001010111100000;
			5'h04: rd_q <= 168'b011110111010110110111000011100110011100010110001100011011100101100000010101001110110001110111010111100111010111101100110110000010101110000000110101110011000010110010100;
			5'h03: rd_q <= 168'b101000001111011000110001111101111100011110000000011111110100110100001001101110110010110010001001001011000010111111010000100111000110100011000001011000110010010110110111;
			5'h02: rd_q <= 168'b111010101110001111111011001101010001001001101001010110001000101011010100110100010000110001110010001001010011111001111100010010110101111101111100100000011000000100010010;
			5'h01: rd_q <= 168'b110000101000101010001001111011000011110110010010100000100001110100100011101000100000010010101000011110111000000001110010000110010010001000101100011001010000010010111010;
			5'h00: rd_q <= 168'b011011010101100001110001100111011011000111100100111101111001100110001011001111000010111000111000010110011010110011100101010110000000100010010011100100110001001001011101;
		default:rd_q <= 168'b0;
		endcase
	end
end

endmodule
