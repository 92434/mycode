
`timescale 1ns / 1ps
module F_short_t12_next_Rom4(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[167:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 168'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h14: rd_q <= 168'b100001101001001010110111001000011010111110100000011100100000110010011010111010110010100011101001110101001010001110111010001010101111111010010111010100000010001111100010;
			5'h13: rd_q <= 168'b111111110011101011001101100100111010111010101010010010010100110001010010101011110111011101000101010110101100100010110101000010000000011011110010100000110110110001011000;
			5'h12: rd_q <= 168'b100100101101100110011110111111010100000101110010001001100110110010000100011110001011111100100110000001111001000110111011001011010011010110111011010110011100100001001110;
			5'h11: rd_q <= 168'b000100111001110101001100001010011111000011001101001011000100000001000000101011010010100100111110100001110011100001110011010100110000011010110000101000011000011000100000;
			5'h10: rd_q <= 168'b100011001101101100100011111001010011100011101110110000000011010001110011110010110001100110011100101000010001000011100110100000001100110000000100100111010011011000000100;
			5'h0f: rd_q <= 168'b010000111100010110000000101100110011001011101000110101111100011001111001000001100101111101101101011101101111000011001101111100111111111110000111101011001000110011000111;
			5'h0e: rd_q <= 168'b011100100111110001100101001111000011101011111110110000110001001100111110111010110011110100001100110010001001101110110100000101110110110011000011000100011011000111111001;
			5'h0d: rd_q <= 168'b111110010011111011100100110101101101010000011000011110000101000010100110110011110000110111100010000000011110010100101010110001111111111111111101100110010010110001101110;
			5'h0c: rd_q <= 168'b100111110011111000010101111110101100101001000110010010110000011001001111000001000010101000111001110111001010100111011001001100010111001101111000110010101101000101000110;
			5'h0b: rd_q <= 168'b100101010000001000011100100000110101100011100110011010100010000110110000100011010111110101000010010011000100000011110001000110111110010001100001001100100011011011011011;
			5'h0a: rd_q <= 168'b111100010001010100010001010001011111101001101011100000000010100000010111011110011101000011101001000101101001100010001100011011011100101010000101000110011101011010010001;
			5'h09: rd_q <= 168'b101000010011011111001000011011111110011010010101011010101010001001111111100000101110000110110001111101101010110001101011111011011110100001100101010011110011001101101000;
			5'h08: rd_q <= 168'b010110000010101101110010000001010010010010101011000100101101101101000000000110111111110001011111101000110110000111101110011110011000000011010110111101010101100001010010;
			5'h07: rd_q <= 168'b100100001110100000001101001000001111100001010111101110001111001000111001001100100010110010111010000011111010010100001011010000000001110001011000001000101101001101100010;
			5'h06: rd_q <= 168'b010110101000110000101111101000100100010000011010010011111100110000111010000001010110101110000101101110100101010111111110001011110111010101000111100101110101100010101010;
			5'h05: rd_q <= 168'b001010111010010000101000011011110111011100010010011110011101100001000011111000000101001100001101101110111010011011011111101011011111000101000101111011100010101111000000;
			5'h04: rd_q <= 168'b111101110101101101110000111001100111000101100011000110111001011000000101010011101100011101110101111001110101111011001101100000101011100000001101011100110000101100101000;
			5'h03: rd_q <= 168'b000010101010110101010010111110000101100011001111000111000000111100111111011001011101001010011011001111101101001100111010000101001110001100101101011100001100011101101011;
			5'h02: rd_q <= 168'b100111101000011011000111011111011111001100011101010100111000000010000101101100011001001101101101001011001111000001100011101110101000110001010110101101011000111000100001;
			5'h01: rd_q <= 168'b110011100101010000100010110011111010110011101010111001101010111101101011010101111000001011011001100100011000110001111111000111100111011011110111011111001000010101110001;
			5'h00: rd_q <= 168'b110110101011000011100011001110110110001111001001111011110011001100010110011110000101110001110000101100110101100111001010101100000001000100100111001001100010010010111010;
		default:rd_q <= 168'b0;
		endcase
	end
end

endmodule
