
`timescale 1ns / 1ps
module F_normal_t8_next_Rom0(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[127:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 128'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h0f: rd_q <= 128'b11010100011001101001111100100000101011101011011000111111100110001011110111101001111001001000111011111010101001001110000000111000;
			5'h0e: rd_q <= 128'b11110110011000011110010001100001101110101000100010100010010010111001011001001101110101101001000011111010000010011010111011010010;
			5'h0d: rd_q <= 128'b00101100001100101000111110110100110111010111101100011000010010010001000110100110101011111111011011001010111011010011111000100111;
			5'h0c: rd_q <= 128'b01000001110100000110101010001000000110110110111100101001101111001011100101000001001010100010010110111011101011111100010001101010;
			5'h0b: rd_q <= 128'b00001110010101100010001111100100000000000100101011010100001011100101010110010000011110001111000011110001111110110111001001000111;
			5'h0a: rd_q <= 128'b00011110110110001110011001111100001101110100010010001000010110101010111110001011100101111001011001111110011011111001101000110100;
			5'h09: rd_q <= 128'b10010111011111010100100010000011101111101101010010011101001101010100010010011010100101111100100000000111101000000111110010110110;
			5'h08: rd_q <= 128'b11001011100011111001111100001001101111110001000101000101111101000011100000001000101010100011111010100001110010000110100011000010;
			5'h07: rd_q <= 128'b00110110100000111011001000101011101000001010100001000110010111011011100110110101110101100001101110111011111000100110001111100110;
			5'h06: rd_q <= 128'b10111011100100011111110110000111010101011000001011100001000100000001100110111100010010111010100111010000011100101100011011000110;
			5'h05: rd_q <= 128'b10001110000001010100100000000000110100101101101001000100010100010111101101100110001110110001011111011100101100000110111001101101;
			5'h04: rd_q <= 128'b01111010011111000000100100001001000011001001110010111100000000010110011101111000101010100100100000110000010100000111110010110111;
			5'h03: rd_q <= 128'b10001111011011000110100011001010000111011101111000110110011100110101101101100011001011000011111100100000101001010000010100010111;
			5'h02: rd_q <= 128'b01101110111001100100000001000011010110111101010011000100100001111011101111001100101010100001010000010011101110000010100001011000;
			5'h01: rd_q <= 128'b10101001111100011000110011100110101001011000101101010000100110101111100011000101011110001011101010100011000110111111101000001000;
			5'h00: rd_q <= 128'b11011001100010010000011101011110010000101111100011010111001100011010110011001111101111111011111010101111101011011011010111000001;
		default:rd_q <= 128'b0;
		endcase
	end
end

endmodule
