
`timescale 1ns / 1ps
module F_normal_t10_next_Rom5(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[159:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 160'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h13: rd_q <= 160'b0111001111000011001101001000001011111100010011011101001000100111010101100101010110011011100001101010101010001010110101110011011000111101000010111110111001000010;
			5'h12: rd_q <= 160'b0111110101000001001101111111101100111100101110001110000100111010011011000000100110010111011100111010111110001001110010110101001111110011001000001010100011001100;
			5'h11: rd_q <= 160'b0101100101001101101011110010001110111111010011000000000010000100111000000000110110110100011000010000100010011010100011101011000101111000010001111110111001101011;
			5'h10: rd_q <= 160'b1010010001110100101010100000001010111010010000100001001011010010010001101011101100011001001001010000100110101111110101011010010001101100111111001110100111011001;
			5'h0f: rd_q <= 160'b0110001101000000110101100011000101110101111011101000100001011100100100111000111110110111011010011111110101101011011010101100110000010000111011110110011011111011;
			5'h0e: rd_q <= 160'b1111000110101001000100100101011011011000111100100110010011011111100001101010000011010111110001111010001000100101100001001101100000111100111010100000000001010010;
			5'h0d: rd_q <= 160'b1010000110000010001101011110110100011000001000100000000111111110010011000101101100110000100010001011010100110010100100001010011110000111011011111010000000100111;
			5'h0c: rd_q <= 160'b0111010000011010010101101001000110110000010100010100111101000001001001101001110011101100000000010110001111101011001011101111111111100110100001111010011101010010;
			5'h0b: rd_q <= 160'b1010000100000111100001101010100111011111010010101010001011010101110100101111101100001100101100110111001111110011010111100000110110100000101101011100110110000000;
			5'h0a: rd_q <= 160'b1000100100000111110110101001101100101001000110111100000101010101000101010011100011100101010110100100101110111111101001110110000110111010100100000001110111001011;
			5'h09: rd_q <= 160'b1000011011001101010101110011000001100010111001010110011111101110011001110111010010101011111000011000110011011111111001011000001001010001111100100001010000101011;
			5'h08: rd_q <= 160'b1110000001111000010001000111010001101001111111011111111001001110110011000100100101101111000100011111010101001101101110101101000010000100010011010000100000100000;
			5'h07: rd_q <= 160'b1010101100101111000100100001111010010100100111000101010011110100011111100001110011010000101011000101011100001010000011001000101010001010011110001100111100001111;
			5'h06: rd_q <= 160'b0011100001011001111110001110100101011011101100111111110001010000101100001101010100000101001011110101010011100011111110010011111111101011011000011110111010111110;
			5'h05: rd_q <= 160'b0101001110110100010000010100100100000011001001000101000100001001001010011101110001100001011011110110000000001110000100001001000000010001111100000110011100001101;
			5'h04: rd_q <= 160'b0000000101000000111110011111101101110010000000101010110101000110111001101010100000001000010111011100001010010001100101101011100011101111011111111001000100110111;
			5'h03: rd_q <= 160'b1010100011111011111111000110110101010110100001010011000010011111010001101011010001001101100011101110110100101111011110010101111001100011101000010101111001100110;
			5'h02: rd_q <= 160'b1010010110010110010100011110101111001111101010100101001011110101101100101001110001110100111000000100101110111011111110001111101111111100100010010110111000111001;
			5'h01: rd_q <= 160'b0000010111111011111011010000001100111100110010000000011100011010101001000011010000011000101110101111101001111100010000011111000101111001001010110110110101111110;
			5'h00: rd_q <= 160'b1001111011111100010100001100111110101001111001011110010011111110010000110101011110010001000011110111000100001010111100010000100010110011110010101101000110001011;
		default:rd_q <= 160'b0;
		endcase
	end
end

endmodule
