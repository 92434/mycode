
`timescale 1ns / 1ps
module F_normal_t8_next_Rom7(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[127:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 128'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h0f: rd_q <= 128'b01000100000011101111011010000010001010000111110100111011101001100101011101001000011001000011110000000001010110101001110111010101;
			5'h0e: rd_q <= 128'b01011000011001010001111101101001101110101111011000110000100100100010001101001101010111111110110110010101110110100111110001001110;
			5'h0d: rd_q <= 128'b10000011101000001101010100010000001101101101111001010011011110010111001010000010010101000100101101110111010111111000100011010100;
			5'h0c: rd_q <= 128'b00011100101011000100011111001000000000001001010110101000010111001010101100100000111100011110000111100011111101101110010010001110;
			5'h0b: rd_q <= 128'b00111101101100011100110011111000011011101000100100010000101101010101111100010111001011110010110011111100110111110011010001101000;
			5'h0a: rd_q <= 128'b10000110001101111010111101000110001000001100010101000101010110111111001011100110111001101000110111111010000010010011100100011101;
			5'h09: rd_q <= 128'b00111111110100100000000001010010001000110100111011110100110110010000101111000010100111010110000010110110110110010001000111110101;
			5'h08: rd_q <= 128'b01101101000001110110010001010111010000010101000010001100101110110111001101101011101011000011011101110111110001001100011111001100;
			5'h07: rd_q <= 128'b11011111111011101100010101001111111101100110100110111101000100010100100010101011010111100100111001010101101011000100110111111101;
			5'h06: rd_q <= 128'b10110100110001111010111001000000111110001101100011110111100100111000110100011111101111110011001001001100001010010001110010101011;
			5'h05: rd_q <= 128'b11110100111110000001001000010010000110010011100101111000000000101100111011110001010101001001000001100000101000001111100101101110;
			5'h04: rd_q <= 128'b10110110000101011110111111010101011001101101000000010011110101111100110100010101100100010110001110110100000000111100101001011111;
			5'h03: rd_q <= 128'b11011101110011001000000010000110101101111010100110001001000011110111011110011001010101000010100000100111011100000101000010110000;
			5'h02: rd_q <= 128'b11111011001011100010011110001100000101100111101011011110000001001000101001011001001110000110100010110011011111100011010001100001;
			5'h01: rd_q <= 128'b00011011110111110011000011111101110110001001110111010001010100100010001001001100101101100110000010101010000100101010101111110011;
			5'h00: rd_q <= 128'b01011101110010000110000000101010010000101100100110111001011110100111000000100000101100111000100110000101010011101000000011111001;		default:rd_q <= 128'b0;
		endcase
	end
end

endmodule
