
`timescale 1ns / 1ps
module F_short_t12_next_Rom6(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[167:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 168'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h14: rd_q <= 168'b100001000000010000110101010000111000000000001111111011011100100110110000101100110000111111111110110001100110111010100011000111001010011011110010000011110100111011111010;
			5'h13: rd_q <= 168'b001111111100111010110011011001001110101110101010100100100101001100010100101010111101110111010001010101101011001000101101010000100000000110111100101000001101101100010110;
			5'h12: rd_q <= 168'b100000010001011011111111001101001011101110111011011110001101000110110111000101111110101000001101001100101010001000100011010111010101010000111001000011010011010000010001;
			5'h11: rd_q <= 168'b000001001110011101010011000010100111110000110011010010110001000000010000001010110100101001001111101000011100111000011100110101001100000110101100001010000110000110001000;
			5'h10: rd_q <= 168'b001000110011011011001000111110010100111000111011101100000000110100011100111100101100011001100111001010000100010000111001101000000011001100000001001001110100110110000001;
			5'h0f: rd_q <= 168'b111001111000000110110100111000101101001010101110001111000001111001000011010011001011000011111101101101110101100101011000001000011110101000011101110111011100011000110010;
			5'h0e: rd_q <= 168'b010011100100111101010101000010101111101101001100010010000110000110000100101111100010110110100001011010111000010111001011110011101101011110011011001010011100111101111111;
			5'h0d: rd_q <= 168'b100110111110111100100001101111100101111011100001111011110101111010111111101110100000011010111100001100110011111100000111001001111110011010101000101111010000110100011001;
			5'h0c: rd_q <= 168'b100000100110111100011101111101010101100101110110011000111000101100000101110010001100111101001010110001000110110000111011110110100100010110001001111010011111001001010011;
			5'h0b: rd_q <= 168'b110100100011000001010011111011101100100000101101100100110110011110110001001011100111100001110110011110011111010101010111000110111110110011100100011110100110100010110101;
			5'h0a: rd_q <= 168'b011011101001010100001000000101001000101101101001000110001010111101001110110110101001011011011000000111000000010100000101110100000111111000001010101010111101011010100101;
			5'h09: rd_q <= 168'b001010000100110111110010000110111111100110100101010110101010100010011111111000001011100001101100011111011010101100011010111110110111101000011001010100111100110011011010;
			5'h08: rd_q <= 168'b101100111010101001000100000010101010001011001101001101011111110001000110000011110011101011010011010110111001111000110110000010000111100101100010011001100001000000010110;
			5'h07: rd_q <= 168'b100000011001101010011011110000111101010111110010000111110111011000011000010001010100111011101010001100001010111100001111010001100001111001000001110100111111001011011010;
			5'h06: rd_q <= 168'b101100110000001110010011011000110111101011100001011000101011100110011000100010001001111100100101110111011101001100110010000111011100010000000110001111101001000000101000;
			5'h05: rd_q <= 168'b000010101110100100001010000110111101110111000100100111100111011000010000111110000001010011000011011011101110100110110111111010110111110001010001011110111000101011110000;
			5'h04: rd_q <= 168'b001111011101011011011100001110011001110001011000110001101110010110000001010100111011000111011101011110011101011110110011011000001010111000000011010111001100001011001010;
			5'h03: rd_q <= 168'b111101011101101110000000011100000000100000100111110011101110110000010010110101000101001110000000001001010101000110100101110110000010110100110111011010101101010011011001;
			5'h02: rd_q <= 168'b011101010111000111111101100110101000100100110100101011000100010101101010011010001000011000111001000100101001111100111110001001011010111110111110010000001100000010001001;
			5'h01: rd_q <= 168'b011000010100010101000100111101100001111011001001010000010000111010010001110100010000001001010100001111011100000000111001000011001001000100010110001100101000001001011101;
			5'h00: rd_q <= 168'b100100110000110010100000010001010011001100010101100010101000011001010011100101111101001011011000100111111001000000111111001110100001110100011110000100101100111100101100;
		default:rd_q <= 168'b0;
		endcase
	end
end

endmodule
