
`timescale 1ns / 1ps
module F_normal_t12_next_Rom1(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b011100111101010100100000001100110111011111010000111100010110000001001000100010000101011000011101100011011001101001111001100001010001110001000101000111010001000011100000101110000011001000111001;
			5'h16: rd_q <= 192'b101001010110111010000111111010011000010010110110111010010001111000010001001011111111011110000100010100101011001010101101011110101100100111001100000010101010001100010000111010101001001011001001;
			5'h15: rd_q <= 192'b100000001010011111100100010110110011100001011001110010111110111001011001000100000110111010101100011011101100011000100111000011011111111100101010010010100111100011101011011010001101010111111011;
			5'h14: rd_q <= 192'b011101100011100100101000010101010100110111110100011000111111001100100001001111111010000011111010011000110111011110100010000100000111110011101101010110100001011101010010110111111111100010010110;
			5'h13: rd_q <= 192'b010000001001000011010110000001100101101101001100111010110000001010010000001100001000111110100001001101000011001000001001100000010101100010110101101001000101100100010010101011111011000000101000;
			5'h12: rd_q <= 192'b000011100011101000110100110100000110100010100001010100101100011100001011100000010011101001001100000100001000011101111101001110010010001011010000000101100000011001000101000001011010100111110111;
			5'h11: rd_q <= 192'b001010010011101010111011101001101000111011101111001111111101100001111011000110101101011010011000110000100101001011010000110001000110111100001010100001101110010010010110101001110011011100100101;
			5'h10: rd_q <= 192'b100101011001100100001110011011101111001100100000101111110101101010000000110000011100000110101000011110000101101010110001101110011111010011010001001110011100001110000110110111000001000110110100;
			5'h0f: rd_q <= 192'b110110011110100000011011011100100000110111000111101101011101100111101011010111001100001110010101101011010101100000110010111000010101111010011000001101000100000101111100101000010010001001011100;
			5'h0e: rd_q <= 192'b010000111010000110101110001101001110011110110010010111110101111110111000101111101010111001110010101101111001000011110101110111011000000101110101111110011101111111000011100001000000111101100011;
			5'h0d: rd_q <= 192'b001011100100101001110010001111110101110100011101001000111100001111100111001000010110110001101101001001000010110001100000110101001101101001101101011100101101101001000001001010100011010110100000;
			5'h0c: rd_q <= 192'b001110011100010011011010011010111000010010110101011001011001001111100111101000110000101001100010101010111110100100010000101000100101101011111000111000111111101010101010000111010011001100101001;
			5'h0b: rd_q <= 192'b110010100000010011111110001011000111011001100001010000011011001010111000001010101001111101000010110000110110100000111001111101111011010111011110111011010000100100100010001101100000100101111111;
			5'h0a: rd_q <= 192'b000111100110111010110001011100111010011111100011100110010101011100100011111111000101110011110000101110111111111101001100011100101000110000110111101001010011010111110101100010110001101111011110;
			5'h09: rd_q <= 192'b111000110001011111010101110101010011000011000101100010011100010011000000111111111001011110110110110111110011101001111000000100100011001100100000011101001011110101111101100010111010110111011011;
			5'h08: rd_q <= 192'b101010000001101001001000000110111001011110110101011001011100000110111110111100101100100000110110101001000011111110010001100001111101010110001001111001001000000000100110011001010110011010000000;
			5'h07: rd_q <= 192'b111001110000001001011010001011101111010000110110010101111010010101010000101011100101111011110011001011011001000011001100100110111011111101011111101100111100010101000001010101100000000100010100;
			5'h06: rd_q <= 192'b111000000111000000010000001111111111011000101000110110111000000100110000110010001000011100000100001100001100000011000100010111101111001011110001001101000100001100001010001110101011000101010000;
			5'h05: rd_q <= 192'b000111000001010100111000000111001110001000000010000101001000001110010011000100101101110100000000011001110101011001011110101001010001100111100011101101100111000001111011001001000011011000111111;
			5'h04: rd_q <= 192'b011011010110110110000000100001101110000010100111000010110110001001011010010111110011001010101111011101001100000100001011100100001100001011011110100001010111111001101100011010100011101111011000;
			5'h03: rd_q <= 192'b001010110000100000010001100100111000111000000110111111011100111101011101001011010110101101111000101110110110110000101100100110001111101001111001101101001110101100101010000010010111100111101110;
			5'h02: rd_q <= 192'b010100100100001000001011001101010010111010000001001110111110100010110111011111111000001000101110011001000011111111000011010111100011010010101010110101000101000111001010111011100110110001100000;
			5'h01: rd_q <= 192'b101011011100011110110010010001110001011010110111111010100010101100010101011010111010111010101010011111100000011110001001100011101111010011011001000000110110110100000000010111101010000100111011;
			5'h00: rd_q <= 192'b111000100110101100101000010101101100100110101011100111100111001000111101111010110010000100011100111100111100100111101001001100011101101100101001100011100110111101100110111111001001100010101001;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
