`timescale 1ns / 1ps
module F_normal_t10_next_Rom1(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[159:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 160'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h13: rd_q <= 160'b0100010011010011011011101000111011000000011000100100010111111011111000000111010100001111001010110111110001100110001010100001111111011011100110000101010000000011;
			5'h12: rd_q <= 160'b1010110011110011010110010001001011001111001100010111010000101000010001011011010111000000011110110010110001010111111011000100001100111001001011000011110011100011;
			5'h11: rd_q <= 160'b1100101010100001101000001110110011110011011011010100000000011111100001100101111110001000000010101011111001010010111000101001010101010011100110101111011010001001;
			5'h10: rd_q <= 160'b1111101110111100000001011000010110101011011110111011110110000111011001101011100000001110011001001111010100001001010010010100001101100000000001101011110111100010;
			5'h0f: rd_q <= 160'b0101111110100000111111111000110101011011110111101111010110101000001111000000001111111101011100111111001111100101010111011100001001101011101100011000111110011110;
			5'h0e: rd_q <= 160'b1111100000011100110100100001010010000111110100011001010100001010111000011000000000101110010101000111101001010110010101110000010010110110100011000011010101101011;
			5'h0d: rd_q <= 160'b1010010011010101111110110111111110001101011110101000111101000111110010001011101010010100101111110011110011011101000110010111110111011001001100100010001000000010;
			5'h0c: rd_q <= 160'b0011100101000101010011111011101000000001101010111001001110011100111011001110001001110111010101111110101001111001101101101000001001100011010111001100010100000011;
			5'h0b: rd_q <= 160'b1010110010001110110011110011001111111011111100001011110111111110001000101011100101010111000000110101000011000001111100111101111110100100100101001111100001110010;
			5'h0a: rd_q <= 160'b0000101000010000011110000110101010011101111101001010101000101101010111010010111110110000110010110011011100111111001101011110000011011010000010110101110011011000;
			5'h09: rd_q <= 160'b1111011010111000101000101101111000100010000111101100000110011010011110011110101101011011011101110100000100111011000110111101111001101100001010111100001011011000;
			5'h08: rd_q <= 160'b1111011001000100000010100000010010010110101000010010101111110001110011101100111110011111100111001111110101001101000111111111000001010010100111011110001001000110;
			5'h07: rd_q <= 160'b0000111000000111100001000100011101000110100111111101111111100100111011001100010010010110111100010001111101010100110110111010110100001000010001001101000010000010;
			5'h06: rd_q <= 160'b1011000001001001010000001101100010111001101001001111110100111011100011110010110000010111000000110101110010010110011010110111111100000100101111010001101111110111;
			5'h05: rd_q <= 160'b0110010100111111010001100100011100110101111010000101100011000011000110110100001011011000111011000011011100011011000000001000001111001000111000100110000011101001;
			5'h04: rd_q <= 160'b0001010000001111100111111011011100100000001010101101010001101110011010101000000010000101110111000010100100011001011010111000111011110111111110010001001101110000;
			5'h03: rd_q <= 160'b0011001101001001011000110111101101100111000010011001100101010111011001100100110101000100110110101011110100000011100001101110001110010101110111011100011000010010;
			5'h02: rd_q <= 160'b1110010110010011101110110001001011110101111111111011111111111000001001001100111011010010001100001101010001001011100111001011101001100111010111101100001111100010;
			5'h01: rd_q <= 160'b0101111110111110110100000011001111001100100000000111000110101010010000110100000110001011101011111010011111000100000111110001011110010010101101101101011111100000;
			5'h00: rd_q <= 160'b0110011011100101011001110001100110010011100111111110011101110111101110100000110011001001001101010110110111110010111110110000111100100001110001101100100011010101;
		default:rd_q <= 160'b0;
		endcase
	end
end

endmodule
