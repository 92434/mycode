
`timescale 1ns / 1ps
module F_normal_t8_next_Rom3(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[127:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 128'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h0f: rd_q <= 128'b00011010100011001101001111100100000101011101011011000111111100110001011110111101001111001001000111011111010101001001110000000111;
			5'h0e: rd_q <= 128'b01110100111111110111001100011100011000000000101000001011100001010010110000111101010010001001010101100010000100110100010111000110;
			5'h0d: rd_q <= 128'b10001110110010100010011010001110010010011110111111001100101110111110111001010011101110100001010011100000000000100000111111101110;
			5'h0c: rd_q <= 128'b01100010000010010100001011000001010101000011011011111010111110111100100111011100110101110000001111001010001001111000100010010001;
			5'h0b: rd_q <= 128'b10001010100001101011001100000100010100100100100111110101001101110000011011010101011000001111010000100111011000001100011001100010;
			5'h0a: rd_q <= 128'b11010111101111011000001111101111001010000101111010101110100100111110100000011000100101100111110000110101011010010001001101111110;
			5'h09: rd_q <= 128'b10101100101110100111100110100000100011100011011110110011111100100100101110001110010001000011000010000111000000101001111110110010;
			5'h08: rd_q <= 128'b01110011010000101011110001110001011000001011100100110111011100101101100111110101111001110000000010101001011010110111110100000100;
			5'h07: rd_q <= 128'b10111000100001011010011011110101100011011111100000101000100111110101010000101011101011000000101011110000100010101101110001011000;
			5'h06: rd_q <= 128'b10101001001001111110111100000000000100110101110101111100011101101110000000101010100111111011110010111101111110001100100011111100;
			5'h05: rd_q <= 128'b11110000101111111001000111101000100111110100000011111000111101001011110111111111010110101100111110111111100110111101010111111011;
			5'h04: rd_q <= 128'b10000100000000111111011001011001111100111101001100111000001100101110000010001000011110101010001100111111010101011010011110111100;
			5'h03: rd_q <= 128'b10011010101000011111101001100001100100011111101101101001011111001010011100001011000010100110110111011101010010110000100010001000;
			5'h02: rd_q <= 128'b00001101110111001100100000001000011010110111101010011000100100001111011101111001100101010100001010000010011101110000010100001011;
			5'h01: rd_q <= 128'b00010101001111100011000110011100110101001011000101101010000100110101111100011000101011110001011101010100011000110111111101000001;
			5'h00: rd_q <= 128'b00101110001010001000011100100011111000111111001010010101000000000001101011100011100011101101010001101011010111001000111010110110;
		default:rd_q <= 128'b0;
		endcase
	end
end

endmodule
