`timescale 1ns / 1ps
module F_normal_t10_next_Rom3(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[159:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 160'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h13: rd_q <= 160'b1101110001000001011010000011000011110000101111100101111101110010110110001000001001010010101101110101101110110011111101001010011110011010010011101110100100000101;
			5'h12: rd_q <= 160'b1110011001001001011001011101011111110011011010101001001100000110001100011111001001100001011000110100111110111111100001010011000010100010111000111111001100111101;
			5'h11: rd_q <= 160'b0111011001111011000001101011010111111100101110010001010111111100000000011110001011101101001010011101001111110010100100101011101010001111011111101110100110100001;
			5'h10: rd_q <= 160'b1011011101001001110111000111110011101010000110100110010010010110000110010100010000011101110011111100010110001110000001100110111101101111001100010000011101111110;
			5'h0f: rd_q <= 160'b1001111001001110111000101111111011010110001100110011011010011101110011111110101011100001000010100000010000110101000000110100111100101101110111001100101111100001;
			5'h0e: rd_q <= 160'b1111001101110010100001110001011001100001010100101010101101001110100110001111111100011010111010001001101000111111111010111110000101000001000010111111000101011111;
			5'h0d: rd_q <= 160'b1010000010010011101000111100001001100011100110100010100000100110001100101100010010111011011110010011011111111011000100100110000011000001011111000010000010000110;
			5'h0c: rd_q <= 160'b1100001100100100111000000111110111000000110011000010101011101011000110111010011110001100101010000111111000110100000100111000000011110100011111111100110101000101;
			5'h0b: rd_q <= 160'b1010001010000101011011101101000101111110001110001010010010001000010010000100010001001011100101100010110011111100001010001100100001011110000101011001011000011010;
			5'h0a: rd_q <= 160'b0000001010000100000111100001101010100111011111010010101010001011010101110100101111101100001100101100110111001111110011010111100000110110100000101101011100110110;
			5'h09: rd_q <= 160'b0011110110101110001010001011011110001000100001111011000001100110100111100111101011010110110111011101000001001110110001101111011110011011000010101111000010110110;
			5'h08: rd_q <= 160'b1011010000110111110111111001110010100101011011001100000100001011101100110101100111111001101100011100011110011111000100111100001110100011100101111101000010010111;
			5'h07: rd_q <= 160'b1000101000100111001111000000110001010001011000110111110000001110111110111101101100111011111010101011111100011001011000101101010011110101001000011001110000100110;
			5'h06: rd_q <= 160'b1110000101100111111000111010010101101110110011111111000101000010110000110101010000010100101111010101001110001111111001001111111110101101100001111011101011111000;
			5'h05: rd_q <= 160'b0101110110011100101111110001111100001101000110000101001111001011001001101010010110111001000100000111000110100000111010100011111100101001101000001100110000111001;
			5'h04: rd_q <= 160'b0000010100000011111001111110110111001000000010101011010100011011100110101010000000100001011101110000101001000110010110101110001110111101111111100100010011011100;
			5'h03: rd_q <= 160'b1000010101110100100001011100001101011001000001101110110110100010000110010111100101001111011000000101011110001100101101011000011101010010010001111101100110000010;
			5'h02: rd_q <= 160'b1011000011000010001100111101100100111101101110110110010000001001110010011101100110101010110110101100110111011110101100110001000100101110111001110001100011111110;
			5'h01: rd_q <= 160'b0001011111101111101101000000110011110011001000000001110001101010100100001101000001100010111010111110100111110001000001111100010111100100101011011011010111111000;
			5'h00: rd_q <= 160'b0101110101101010001101110100100010100100100001011011110000100110000011101111011000111101011001100010011100011010100101001101110000010011111010011110011000110110;
		default:rd_q <= 160'b0;
		endcase
	end
end

endmodule
