`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2016/01/01 09:04:08
// Design Name: 
// Module Name: ldpc_check_ram_v
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ldpc_check_ram_noip(
    input aclr,
    input clock,
    input [44:0] data,
    input [7:0] rdaddress,
    input rden,
    input [7:0] wraddress,
    input wren,
    output reg [44:0] q
    );
    
    reg [44:0] ram_buff_00;
    reg [44:0] ram_buff_01;
    reg [44:0] ram_buff_02;
    reg [44:0] ram_buff_03;
    reg [44:0] ram_buff_04;
    reg [44:0] ram_buff_05;
    reg [44:0] ram_buff_06;
    reg [44:0] ram_buff_07;
    reg [44:0] ram_buff_08;
    reg [44:0] ram_buff_09;
    reg [44:0] ram_buff_0A;
    reg [44:0] ram_buff_0B;
    reg [44:0] ram_buff_0C;
    reg [44:0] ram_buff_0D;
    reg [44:0] ram_buff_0E;
    reg [44:0] ram_buff_0F;
    reg [44:0] ram_buff_10;
    reg [44:0] ram_buff_11;
    reg [44:0] ram_buff_12;
    reg [44:0] ram_buff_13;
    reg [44:0] ram_buff_14;
    reg [44:0] ram_buff_15;
    reg [44:0] ram_buff_16;
    reg [44:0] ram_buff_17;
    reg [44:0] ram_buff_18;
    reg [44:0] ram_buff_19;
    reg [44:0] ram_buff_1A;
    reg [44:0] ram_buff_1B;
    reg [44:0] ram_buff_1C;
    reg [44:0] ram_buff_1D;
    reg [44:0] ram_buff_1E;
    reg [44:0] ram_buff_1F;
    reg [44:0] ram_buff_20;
    reg [44:0] ram_buff_21;
    reg [44:0] ram_buff_22;
    reg [44:0] ram_buff_23;
    reg [44:0] ram_buff_24;
    reg [44:0] ram_buff_25;
    reg [44:0] ram_buff_26;
    reg [44:0] ram_buff_27;
    reg [44:0] ram_buff_28;
    reg [44:0] ram_buff_29;
    reg [44:0] ram_buff_2A;
    reg [44:0] ram_buff_2B;
    reg [44:0] ram_buff_2C;
    reg [44:0] ram_buff_2D;
    reg [44:0] ram_buff_2E;
    reg [44:0] ram_buff_2F;
    reg [44:0] ram_buff_30;
    reg [44:0] ram_buff_31;
    reg [44:0] ram_buff_32;
    reg [44:0] ram_buff_33;
    reg [44:0] ram_buff_34;
    reg [44:0] ram_buff_35;
    reg [44:0] ram_buff_36;
    reg [44:0] ram_buff_37;
    reg [44:0] ram_buff_38;
    reg [44:0] ram_buff_39;
    reg [44:0] ram_buff_3A;
    reg [44:0] ram_buff_3B;
    reg [44:0] ram_buff_3C;
    reg [44:0] ram_buff_3D;
    reg [44:0] ram_buff_3E;
    reg [44:0] ram_buff_3F;
    reg [44:0] ram_buff_40;
    reg [44:0] ram_buff_41;
    reg [44:0] ram_buff_42;
    reg [44:0] ram_buff_43;
    reg [44:0] ram_buff_44;
    reg [44:0] ram_buff_45;
    reg [44:0] ram_buff_46;
    reg [44:0] ram_buff_47;
    reg [44:0] ram_buff_48;
    reg [44:0] ram_buff_49;
    reg [44:0] ram_buff_4A;
    reg [44:0] ram_buff_4B;
    reg [44:0] ram_buff_4C;
    reg [44:0] ram_buff_4D;
    reg [44:0] ram_buff_4E;
    reg [44:0] ram_buff_4F;
    reg [44:0] ram_buff_50;
    reg [44:0] ram_buff_51;
    reg [44:0] ram_buff_52;
    reg [44:0] ram_buff_53;
    reg [44:0] ram_buff_54;
    reg [44:0] ram_buff_55;
    reg [44:0] ram_buff_56;
    reg [44:0] ram_buff_57;
    reg [44:0] ram_buff_58;
    reg [44:0] ram_buff_59;
    reg [44:0] ram_buff_5A;
    reg [44:0] ram_buff_5B;
    reg [44:0] ram_buff_5C;
    reg [44:0] ram_buff_5D;
    reg [44:0] ram_buff_5E;
    reg [44:0] ram_buff_5F;
    reg [44:0] ram_buff_60;
    reg [44:0] ram_buff_61;
    reg [44:0] ram_buff_62;
    reg [44:0] ram_buff_63;
    reg [44:0] ram_buff_64;
    reg [44:0] ram_buff_65;
    reg [44:0] ram_buff_66;
    reg [44:0] ram_buff_67;
    reg [44:0] ram_buff_68;
    reg [44:0] ram_buff_69;
    reg [44:0] ram_buff_6A;
    reg [44:0] ram_buff_6B;
    reg [44:0] ram_buff_6C;
    reg [44:0] ram_buff_6D;
    reg [44:0] ram_buff_6E;
    reg [44:0] ram_buff_6F;
    reg [44:0] ram_buff_70;
    reg [44:0] ram_buff_71;
    reg [44:0] ram_buff_72;
    reg [44:0] ram_buff_73;
    reg [44:0] ram_buff_74;
    reg [44:0] ram_buff_75;
    reg [44:0] ram_buff_76;
    reg [44:0] ram_buff_77;
    reg [44:0] ram_buff_78;
    reg [44:0] ram_buff_79;
    reg [44:0] ram_buff_7A;
    reg [44:0] ram_buff_7B;
    reg [44:0] ram_buff_7C;
    reg [44:0] ram_buff_7D;
    reg [44:0] ram_buff_7E;
    reg [44:0] ram_buff_7F;
    reg [44:0] ram_buff_80;
    reg [44:0] ram_buff_81;
    reg [44:0] ram_buff_82;
    reg [44:0] ram_buff_83;
    reg [44:0] ram_buff_84;
    reg [44:0] ram_buff_85;
    reg [44:0] ram_buff_86;
    reg [44:0] ram_buff_87;
    reg [44:0] ram_buff_88;
    reg [44:0] ram_buff_89;
    reg [44:0] ram_buff_8A;
    reg [44:0] ram_buff_8B;
    reg [44:0] ram_buff_8C;
    reg [44:0] ram_buff_8D;
    reg [44:0] ram_buff_8E;
    reg [44:0] ram_buff_8F;
    reg [44:0] ram_buff_90;
    reg [44:0] ram_buff_91;
    reg [44:0] ram_buff_92;
    reg [44:0] ram_buff_93;
    reg [44:0] ram_buff_94;
    reg [44:0] ram_buff_95;
    reg [44:0] ram_buff_96;
    reg [44:0] ram_buff_97;
    reg [44:0] ram_buff_98;
    reg [44:0] ram_buff_99;
    reg [44:0] ram_buff_9A;
    reg [44:0] ram_buff_9B;
    reg [44:0] ram_buff_9C;
    reg [44:0] ram_buff_9D;
    reg [44:0] ram_buff_9E;
    reg [44:0] ram_buff_9F;
    reg [44:0] ram_buff_A0;
    reg [44:0] ram_buff_A1;
    reg [44:0] ram_buff_A2;
    reg [44:0] ram_buff_A3;
    reg [44:0] ram_buff_A4;
    reg [44:0] ram_buff_A5;
    reg [44:0] ram_buff_A6;
    reg [44:0] ram_buff_A7;
    reg [44:0] ram_buff_A8;
    reg [44:0] ram_buff_A9;
    reg [44:0] ram_buff_AA;
    reg [44:0] ram_buff_AB;
    reg [44:0] ram_buff_AC;
    reg [44:0] ram_buff_AD;
    reg [44:0] ram_buff_AE;
    reg [44:0] ram_buff_AF;
    reg [44:0] ram_buff_B0;
    reg [44:0] ram_buff_B1;
    reg [44:0] ram_buff_B2;
    reg [44:0] ram_buff_B3;
    reg [44:0] ram_buff_B4;
    reg [44:0] ram_buff_B5;
    reg [44:0] ram_buff_B6;
    reg [44:0] ram_buff_B7;
    reg [44:0] ram_buff_B8;
    reg [44:0] ram_buff_B9;
    reg [44:0] ram_buff_BA;
    reg [44:0] ram_buff_BB;
    reg [44:0] ram_buff_BC;
    reg [44:0] ram_buff_BD;
    reg [44:0] ram_buff_BE;
    reg [44:0] ram_buff_BF;
    reg [44:0] ram_buff_C0;
    reg [44:0] ram_buff_C1;
    reg [44:0] ram_buff_C2;
    reg [44:0] ram_buff_C3;
    reg [44:0] ram_buff_C4;
    reg [44:0] ram_buff_C5;
    reg [44:0] ram_buff_C6;
    reg [44:0] ram_buff_C7;
    reg [44:0] ram_buff_C8;
    reg [44:0] ram_buff_C9;
    reg [44:0] ram_buff_CA;
    reg [44:0] ram_buff_CB;
    reg [44:0] ram_buff_CC;
    reg [44:0] ram_buff_CD;
    reg [44:0] ram_buff_CE;
    reg [44:0] ram_buff_CF;
    reg [44:0] ram_buff_D0;
    reg [44:0] ram_buff_D1;
    reg [44:0] ram_buff_D2;
    reg [44:0] ram_buff_D3;
    reg [44:0] ram_buff_D4;
    reg [44:0] ram_buff_D5;
    reg [44:0] ram_buff_D6;
    reg [44:0] ram_buff_D7;
    reg [44:0] ram_buff_D8;
    reg [44:0] ram_buff_D9;
    reg [44:0] ram_buff_DA;
    reg [44:0] ram_buff_DB;
    reg [44:0] ram_buff_DC;
    reg [44:0] ram_buff_DD;
    reg [44:0] ram_buff_DE;
    reg [44:0] ram_buff_DF;
    reg [44:0] ram_buff_E0;
    reg [44:0] ram_buff_E1;
    reg [44:0] ram_buff_E2;
    reg [44:0] ram_buff_E3;
    reg [44:0] ram_buff_E4;
    reg [44:0] ram_buff_E5;
    reg [44:0] ram_buff_E6;
    reg [44:0] ram_buff_E7;
    reg [44:0] ram_buff_E8;
    reg [44:0] ram_buff_E9;
    reg [44:0] ram_buff_EA;
    reg [44:0] ram_buff_EB;
    reg [44:0] ram_buff_EC;
    reg [44:0] ram_buff_ED;
    reg [44:0] ram_buff_EE;
    reg [44:0] ram_buff_EF;
    reg [44:0] ram_buff_F0;
    reg [44:0] ram_buff_F1;
    reg [44:0] ram_buff_F2;
    reg [44:0] ram_buff_F3;
    reg [44:0] ram_buff_F4;
    reg [44:0] ram_buff_F5;
    reg [44:0] ram_buff_F6;
    reg [44:0] ram_buff_F7;
    reg [44:0] ram_buff_F8;
    reg [44:0] ram_buff_F9;
    reg [44:0] ram_buff_FA;
    reg [44:0] ram_buff_FB;
    reg [44:0] ram_buff_FC;
    reg [44:0] ram_buff_FD;
    reg [44:0] ram_buff_FE;
    reg [44:0] ram_buff_FF;


    
 always @(posedge clock)begin
        if(aclr)begin
        ram_buff_00 <= 45'h000000000000;
        ram_buff_01 <= 45'h000000000000;
        ram_buff_02 <= 45'h000000000000;
        ram_buff_03 <= 45'h000000000000;
        ram_buff_04 <= 45'h000000000000;
        ram_buff_05 <= 45'h000000000000;
        ram_buff_06 <= 45'h000000000000;
        ram_buff_07 <= 45'h000000000000;
        ram_buff_08 <= 45'h000000000000;
        ram_buff_09 <= 45'h000000000000;
        ram_buff_0A <= 45'h000000000000;
        ram_buff_0B <= 45'h000000000000;
        ram_buff_0C <= 45'h000000000000;
        ram_buff_0D <= 45'h000000000000;
        ram_buff_0E <= 45'h000000000000;
        ram_buff_0F <= 45'h000000000000;
        ram_buff_10 <= 45'h000000000000;
        ram_buff_11 <= 45'h000000000000;
        ram_buff_12 <= 45'h000000000000;
        ram_buff_13 <= 45'h000000000000;
        ram_buff_14 <= 45'h000000000000;
        ram_buff_15 <= 45'h000000000000;
        ram_buff_16 <= 45'h000000000000;
        ram_buff_17 <= 45'h000000000000;
        ram_buff_18 <= 45'h000000000000;
        ram_buff_19 <= 45'h000000000000;
        ram_buff_1A <= 45'h000000000000;
        ram_buff_1B <= 45'h000000000000;
        ram_buff_1C <= 45'h000000000000;
        ram_buff_1D <= 45'h000000000000;
        ram_buff_1E <= 45'h000000000000;
        ram_buff_1F <= 45'h000000000000;
        ram_buff_20 <= 45'h000000000000;
        ram_buff_21 <= 45'h000000000000;
        ram_buff_22 <= 45'h000000000000;
        ram_buff_23 <= 45'h000000000000;
        ram_buff_24 <= 45'h000000000000;
        ram_buff_25 <= 45'h000000000000;
        ram_buff_26 <= 45'h000000000000;
        ram_buff_27 <= 45'h000000000000;
        ram_buff_28 <= 45'h000000000000;
        ram_buff_29 <= 45'h000000000000;
        ram_buff_2A <= 45'h000000000000;
        ram_buff_2B <= 45'h000000000000;
        ram_buff_2C <= 45'h000000000000;
        ram_buff_2D <= 45'h000000000000;
        ram_buff_2E <= 45'h000000000000;
        ram_buff_2F <= 45'h000000000000;
        ram_buff_30 <= 45'h000000000000;
        ram_buff_31 <= 45'h000000000000;
        ram_buff_32 <= 45'h000000000000;
        ram_buff_33 <= 45'h000000000000;
        ram_buff_34 <= 45'h000000000000;
        ram_buff_35 <= 45'h000000000000;
        ram_buff_36 <= 45'h000000000000;
        ram_buff_37 <= 45'h000000000000;
        ram_buff_38 <= 45'h000000000000;
        ram_buff_39 <= 45'h000000000000;
        ram_buff_3A <= 45'h000000000000;
        ram_buff_3B <= 45'h000000000000;
        ram_buff_3C <= 45'h000000000000;
        ram_buff_3D <= 45'h000000000000;
        ram_buff_3E <= 45'h000000000000;
        ram_buff_3F <= 45'h000000000000;
        ram_buff_40 <= 45'h000000000000;
        ram_buff_41 <= 45'h000000000000;
        ram_buff_42 <= 45'h000000000000;
        ram_buff_43 <= 45'h000000000000;
        ram_buff_44 <= 45'h000000000000;
        ram_buff_45 <= 45'h000000000000;
        ram_buff_46 <= 45'h000000000000;
        ram_buff_47 <= 45'h000000000000;
        ram_buff_48 <= 45'h000000000000;
        ram_buff_49 <= 45'h000000000000;
        ram_buff_4A <= 45'h000000000000;
        ram_buff_4B <= 45'h000000000000;
        ram_buff_4C <= 45'h000000000000;
        ram_buff_4D <= 45'h000000000000;
        ram_buff_4E <= 45'h000000000000;
        ram_buff_4F <= 45'h000000000000;
        ram_buff_50 <= 45'h000000000000;
        ram_buff_51 <= 45'h000000000000;
        ram_buff_52 <= 45'h000000000000;
        ram_buff_53 <= 45'h000000000000;
        ram_buff_54 <= 45'h000000000000;
        ram_buff_55 <= 45'h000000000000;
        ram_buff_56 <= 45'h000000000000;
        ram_buff_57 <= 45'h000000000000;
        ram_buff_58 <= 45'h000000000000;
        ram_buff_59 <= 45'h000000000000;
        ram_buff_5A <= 45'h000000000000;
        ram_buff_5B <= 45'h000000000000;
        ram_buff_5C <= 45'h000000000000;
        ram_buff_5D <= 45'h000000000000;
        ram_buff_5E <= 45'h000000000000;
        ram_buff_5F <= 45'h000000000000;
        ram_buff_60 <= 45'h000000000000;
        ram_buff_61 <= 45'h000000000000;
        ram_buff_62 <= 45'h000000000000;
        ram_buff_63 <= 45'h000000000000;
        ram_buff_64 <= 45'h000000000000;
        ram_buff_65 <= 45'h000000000000;
        ram_buff_66 <= 45'h000000000000;
        ram_buff_67 <= 45'h000000000000;
        ram_buff_68 <= 45'h000000000000;
        ram_buff_69 <= 45'h000000000000;
        ram_buff_6A <= 45'h000000000000;
        ram_buff_6B <= 45'h000000000000;
        ram_buff_6C <= 45'h000000000000;
        ram_buff_6D <= 45'h000000000000;
        ram_buff_6E <= 45'h000000000000;
        ram_buff_6F <= 45'h000000000000;
        ram_buff_70 <= 45'h000000000000;
        ram_buff_71 <= 45'h000000000000;
        ram_buff_72 <= 45'h000000000000;
        ram_buff_73 <= 45'h000000000000;
        ram_buff_74 <= 45'h000000000000;
        ram_buff_75 <= 45'h000000000000;
        ram_buff_76 <= 45'h000000000000;
        ram_buff_77 <= 45'h000000000000;
        ram_buff_78 <= 45'h000000000000;
        ram_buff_79 <= 45'h000000000000;
        ram_buff_7A <= 45'h000000000000;
        ram_buff_7B <= 45'h000000000000;
        ram_buff_7C <= 45'h000000000000;
        ram_buff_7D <= 45'h000000000000;
        ram_buff_7E <= 45'h000000000000;
        ram_buff_7F <= 45'h000000000000;
        ram_buff_80 <= 45'h000000000000;
        ram_buff_81 <= 45'h000000000000;
        ram_buff_82 <= 45'h000000000000;
        ram_buff_83 <= 45'h000000000000;
        ram_buff_84 <= 45'h000000000000;
        ram_buff_85 <= 45'h000000000000;
        ram_buff_86 <= 45'h000000000000;
        ram_buff_87 <= 45'h000000000000;
        ram_buff_88 <= 45'h000000000000;
        ram_buff_89 <= 45'h000000000000;
        ram_buff_8A <= 45'h000000000000;
        ram_buff_8B <= 45'h000000000000;
        ram_buff_8C <= 45'h000000000000;
        ram_buff_8D <= 45'h000000000000;
        ram_buff_8E <= 45'h000000000000;
        ram_buff_8F <= 45'h000000000000;
        ram_buff_90 <= 45'h000000000000;
        ram_buff_91 <= 45'h000000000000;
        ram_buff_92 <= 45'h000000000000;
        ram_buff_93 <= 45'h000000000000;
        ram_buff_94 <= 45'h000000000000;
        ram_buff_95 <= 45'h000000000000;
        ram_buff_96 <= 45'h000000000000;
        ram_buff_97 <= 45'h000000000000;
        ram_buff_98 <= 45'h000000000000;
        ram_buff_99 <= 45'h000000000000;
        ram_buff_9A <= 45'h000000000000;
        ram_buff_9B <= 45'h000000000000;
        ram_buff_9C <= 45'h000000000000;
        ram_buff_9D <= 45'h000000000000;
        ram_buff_9E <= 45'h000000000000;
        ram_buff_9F <= 45'h000000000000;
        ram_buff_A0 <= 45'h000000000000;
        ram_buff_A1 <= 45'h000000000000;
        ram_buff_A2 <= 45'h000000000000;
        ram_buff_A3 <= 45'h000000000000;
        ram_buff_A4 <= 45'h000000000000;
        ram_buff_A5 <= 45'h000000000000;
        ram_buff_A6 <= 45'h000000000000;
        ram_buff_A7 <= 45'h000000000000;
        ram_buff_A8 <= 45'h000000000000;
        ram_buff_A9 <= 45'h000000000000;
        ram_buff_AA <= 45'h000000000000;
        ram_buff_AB <= 45'h000000000000;
        ram_buff_AC <= 45'h000000000000;
        ram_buff_AD <= 45'h000000000000;
        ram_buff_AE <= 45'h000000000000;
        ram_buff_AF <= 45'h000000000000;
        ram_buff_B0 <= 45'h000000000000;
        ram_buff_B1 <= 45'h000000000000;
        ram_buff_B2 <= 45'h000000000000;
        ram_buff_B3 <= 45'h000000000000;
        ram_buff_B4 <= 45'h000000000000;
        ram_buff_B5 <= 45'h000000000000;
        ram_buff_B6 <= 45'h000000000000;
        ram_buff_B7 <= 45'h000000000000;
        ram_buff_B8 <= 45'h000000000000;
        ram_buff_B9 <= 45'h000000000000;
        ram_buff_BA <= 45'h000000000000;
        ram_buff_BB <= 45'h000000000000;
        ram_buff_BC <= 45'h000000000000;
        ram_buff_BD <= 45'h000000000000;
        ram_buff_BE <= 45'h000000000000;
        ram_buff_BF <= 45'h000000000000;
        ram_buff_C0 <= 45'h000000000000;
        ram_buff_C1 <= 45'h000000000000;
        ram_buff_C2 <= 45'h000000000000;
        ram_buff_C3 <= 45'h000000000000;
        ram_buff_C4 <= 45'h000000000000;
        ram_buff_C5 <= 45'h000000000000;
        ram_buff_C6 <= 45'h000000000000;
        ram_buff_C7 <= 45'h000000000000;
        ram_buff_C8 <= 45'h000000000000;
        ram_buff_C9 <= 45'h000000000000;
        ram_buff_CA <= 45'h000000000000;
        ram_buff_CB <= 45'h000000000000;
        ram_buff_CC <= 45'h000000000000;
        ram_buff_CD <= 45'h000000000000;
        ram_buff_CE <= 45'h000000000000;
        ram_buff_CF <= 45'h000000000000;
        ram_buff_D0 <= 45'h000000000000;
        ram_buff_D1 <= 45'h000000000000;
        ram_buff_D2 <= 45'h000000000000;
        ram_buff_D3 <= 45'h000000000000;
        ram_buff_D4 <= 45'h000000000000;
        ram_buff_D5 <= 45'h000000000000;
        ram_buff_D6 <= 45'h000000000000;
        ram_buff_D7 <= 45'h000000000000;
        ram_buff_D8 <= 45'h000000000000;
        ram_buff_D9 <= 45'h000000000000;
        ram_buff_DA <= 45'h000000000000;
        ram_buff_DB <= 45'h000000000000;
        ram_buff_DC <= 45'h000000000000;
        ram_buff_DD <= 45'h000000000000;
        ram_buff_DE <= 45'h000000000000;
        ram_buff_DF <= 45'h000000000000;
        ram_buff_E0 <= 45'h000000000000;
        ram_buff_E1 <= 45'h000000000000;
        ram_buff_E2 <= 45'h000000000000;
        ram_buff_E3 <= 45'h000000000000;
        ram_buff_E4 <= 45'h000000000000;
        ram_buff_E5 <= 45'h000000000000;
        ram_buff_E6 <= 45'h000000000000;
        ram_buff_E7 <= 45'h000000000000;
        ram_buff_E8 <= 45'h000000000000;
        ram_buff_E9 <= 45'h000000000000;
        ram_buff_EA <= 45'h000000000000;
        ram_buff_EB <= 45'h000000000000;
        ram_buff_EC <= 45'h000000000000;
        ram_buff_ED <= 45'h000000000000;
        ram_buff_EE <= 45'h000000000000;
        ram_buff_EF <= 45'h000000000000;
        ram_buff_F0 <= 45'h000000000000;
        ram_buff_F1 <= 45'h000000000000;
        ram_buff_F2 <= 45'h000000000000;
        ram_buff_F3 <= 45'h000000000000;
        ram_buff_F4 <= 45'h000000000000;
        ram_buff_F5 <= 45'h000000000000;
        ram_buff_F6 <= 45'h000000000000;
        ram_buff_F7 <= 45'h000000000000;
        ram_buff_F8 <= 45'h000000000000;
        ram_buff_F9 <= 45'h000000000000;
        ram_buff_FA <= 45'h000000000000;
        ram_buff_FB <= 45'h000000000000;
        ram_buff_FC <= 45'h000000000000;
        ram_buff_FD <= 45'h000000000000;
        ram_buff_FE <= 45'h000000000000;
        ram_buff_FF <= 45'h000000000000;
        end
        else if(wren)begin
            case(wraddress)
            8'h00: ram_buff_00 <= data;
            8'h01: ram_buff_01 <= data;
            8'h02: ram_buff_02 <= data;
            8'h03: ram_buff_03 <= data;
            8'h04: ram_buff_04 <= data;
            8'h05: ram_buff_05 <= data;
            8'h06: ram_buff_06 <= data;
            8'h07: ram_buff_07 <= data;
            8'h08: ram_buff_08 <= data;
            8'h09: ram_buff_09 <= data;
            8'h0A: ram_buff_0A <= data;
            8'h0B: ram_buff_0B <= data;
            8'h0C: ram_buff_0C <= data;
            8'h0D: ram_buff_0D <= data;
            8'h0E: ram_buff_0E <= data;
            8'h0F: ram_buff_0F <= data;
            8'h10: ram_buff_10 <= data;
            8'h11: ram_buff_11 <= data;
            8'h12: ram_buff_12 <= data;
            8'h13: ram_buff_13 <= data;
            8'h14: ram_buff_14 <= data;
            8'h15: ram_buff_15 <= data;
            8'h16: ram_buff_16 <= data;
            8'h17: ram_buff_17 <= data;
            8'h18: ram_buff_18 <= data;
            8'h19: ram_buff_19 <= data;
            8'h1A: ram_buff_1A <= data;
            8'h1B: ram_buff_1B <= data;
            8'h1C: ram_buff_1C <= data;
            8'h1D: ram_buff_1D <= data;
            8'h1E: ram_buff_1E <= data;
            8'h1F: ram_buff_1F <= data;
            8'h20: ram_buff_20 <= data;
            8'h21: ram_buff_21 <= data;
            8'h22: ram_buff_22 <= data;
            8'h23: ram_buff_23 <= data;
            8'h24: ram_buff_24 <= data;
            8'h25: ram_buff_25 <= data;
            8'h26: ram_buff_26 <= data;
            8'h27: ram_buff_27 <= data;
            8'h28: ram_buff_28 <= data;
            8'h29: ram_buff_29 <= data;
            8'h2A: ram_buff_2A <= data;
            8'h2B: ram_buff_2B <= data;
            8'h2C: ram_buff_2C <= data;
            8'h2D: ram_buff_2D <= data;
            8'h2E: ram_buff_2E <= data;
            8'h2F: ram_buff_2F <= data;
            8'h30: ram_buff_30 <= data;
            8'h31: ram_buff_31 <= data;
            8'h32: ram_buff_32 <= data;
            8'h33: ram_buff_33 <= data;
            8'h34: ram_buff_34 <= data;
            8'h35: ram_buff_35 <= data;
            8'h36: ram_buff_36 <= data;
            8'h37: ram_buff_37 <= data;
            8'h38: ram_buff_38 <= data;
            8'h39: ram_buff_39 <= data;
            8'h3A: ram_buff_3A <= data;
            8'h3B: ram_buff_3B <= data;
            8'h3C: ram_buff_3C <= data;
            8'h3D: ram_buff_3D <= data;
            8'h3E: ram_buff_3E <= data;
            8'h3F: ram_buff_3F <= data;
            8'h40: ram_buff_40 <= data;
            8'h41: ram_buff_41 <= data;
            8'h42: ram_buff_42 <= data;
            8'h43: ram_buff_43 <= data;
            8'h44: ram_buff_44 <= data;
            8'h45: ram_buff_45 <= data;
            8'h46: ram_buff_46 <= data;
            8'h47: ram_buff_47 <= data;
            8'h48: ram_buff_48 <= data;
            8'h49: ram_buff_49 <= data;
            8'h4A: ram_buff_4A <= data;
            8'h4B: ram_buff_4B <= data;
            8'h4C: ram_buff_4C <= data;
            8'h4D: ram_buff_4D <= data;
            8'h4E: ram_buff_4E <= data;
            8'h4F: ram_buff_4F <= data;
            8'h50: ram_buff_50 <= data;
            8'h51: ram_buff_51 <= data;
            8'h52: ram_buff_52 <= data;
            8'h53: ram_buff_53 <= data;
            8'h54: ram_buff_54 <= data;
            8'h55: ram_buff_55 <= data;
            8'h56: ram_buff_56 <= data;
            8'h57: ram_buff_57 <= data;
            8'h58: ram_buff_58 <= data;
            8'h59: ram_buff_59 <= data;
            8'h5A: ram_buff_5A <= data;
            8'h5B: ram_buff_5B <= data;
            8'h5C: ram_buff_5C <= data;
            8'h5D: ram_buff_5D <= data;
            8'h5E: ram_buff_5E <= data;
            8'h5F: ram_buff_5F <= data;
            8'h60: ram_buff_60 <= data;
            8'h61: ram_buff_61 <= data;
            8'h62: ram_buff_62 <= data;
            8'h63: ram_buff_63 <= data;
            8'h64: ram_buff_64 <= data;
            8'h65: ram_buff_65 <= data;
            8'h66: ram_buff_66 <= data;
            8'h67: ram_buff_67 <= data;
            8'h68: ram_buff_68 <= data;
            8'h69: ram_buff_69 <= data;
            8'h6A: ram_buff_6A <= data;
            8'h6B: ram_buff_6B <= data;
            8'h6C: ram_buff_6C <= data;
            8'h6D: ram_buff_6D <= data;
            8'h6E: ram_buff_6E <= data;
            8'h6F: ram_buff_6F <= data;
            8'h70: ram_buff_70 <= data;
            8'h71: ram_buff_71 <= data;
            8'h72: ram_buff_72 <= data;
            8'h73: ram_buff_73 <= data;
            8'h74: ram_buff_74 <= data;
            8'h75: ram_buff_75 <= data;
            8'h76: ram_buff_76 <= data;
            8'h77: ram_buff_77 <= data;
            8'h78: ram_buff_78 <= data;
            8'h79: ram_buff_79 <= data;
            8'h7A: ram_buff_7A <= data;
            8'h7B: ram_buff_7B <= data;
            8'h7C: ram_buff_7C <= data;
            8'h7D: ram_buff_7D <= data;
            8'h7E: ram_buff_7E <= data;
            8'h7F: ram_buff_7F <= data;
            8'h80: ram_buff_80 <= data;
            8'h81: ram_buff_81 <= data;
            8'h82: ram_buff_82 <= data;
            8'h83: ram_buff_83 <= data;
            8'h84: ram_buff_84 <= data;
            8'h85: ram_buff_85 <= data;
            8'h86: ram_buff_86 <= data;
            8'h87: ram_buff_87 <= data;
            8'h88: ram_buff_88 <= data;
            8'h89: ram_buff_89 <= data;
            8'h8A: ram_buff_8A <= data;
            8'h8B: ram_buff_8B <= data;
            8'h8C: ram_buff_8C <= data;
            8'h8D: ram_buff_8D <= data;
            8'h8E: ram_buff_8E <= data;
            8'h8F: ram_buff_8F <= data;
            8'h90: ram_buff_90 <= data;
            8'h91: ram_buff_91 <= data;
            8'h92: ram_buff_92 <= data;
            8'h93: ram_buff_93 <= data;
            8'h94: ram_buff_94 <= data;
            8'h95: ram_buff_95 <= data;
            8'h96: ram_buff_96 <= data;
            8'h97: ram_buff_97 <= data;
            8'h98: ram_buff_98 <= data;
            8'h99: ram_buff_99 <= data;
            8'h9A: ram_buff_9A <= data;
            8'h9B: ram_buff_9B <= data;
            8'h9C: ram_buff_9C <= data;
            8'h9D: ram_buff_9D <= data;
            8'h9E: ram_buff_9E <= data;
            8'h9F: ram_buff_9F <= data;
            8'hA0: ram_buff_A0 <= data;
            8'hA1: ram_buff_A1 <= data;
            8'hA2: ram_buff_A2 <= data;
            8'hA3: ram_buff_A3 <= data;
            8'hA4: ram_buff_A4 <= data;
            8'hA5: ram_buff_A5 <= data;
            8'hA6: ram_buff_A6 <= data;
            8'hA7: ram_buff_A7 <= data;
            8'hA8: ram_buff_A8 <= data;
            8'hA9: ram_buff_A9 <= data;
            8'hAA: ram_buff_AA <= data;
            8'hAB: ram_buff_AB <= data;
            8'hAC: ram_buff_AC <= data;
            8'hAD: ram_buff_AD <= data;
            8'hAE: ram_buff_AE <= data;
            8'hAF: ram_buff_AF <= data;
            8'hB0: ram_buff_B0 <= data;
            8'hB1: ram_buff_B1 <= data;
            8'hB2: ram_buff_B2 <= data;
            8'hB3: ram_buff_B3 <= data;
            8'hB4: ram_buff_B4 <= data;
            8'hB5: ram_buff_B5 <= data;
            8'hB6: ram_buff_B6 <= data;
            8'hB7: ram_buff_B7 <= data;
            8'hB8: ram_buff_B8 <= data;
            8'hB9: ram_buff_B9 <= data;
            8'hBA: ram_buff_BA <= data;
            8'hBB: ram_buff_BB <= data;
            8'hBC: ram_buff_BC <= data;
            8'hBD: ram_buff_BD <= data;
            8'hBE: ram_buff_BE <= data;
            8'hBF: ram_buff_BF <= data;
            8'hC0: ram_buff_C0 <= data;
            8'hC1: ram_buff_C1 <= data;
            8'hC2: ram_buff_C2 <= data;
            8'hC3: ram_buff_C3 <= data;
            8'hC4: ram_buff_C4 <= data;
            8'hC5: ram_buff_C5 <= data;
            8'hC6: ram_buff_C6 <= data;
            8'hC7: ram_buff_C7 <= data;
            8'hC8: ram_buff_C8 <= data;
            8'hC9: ram_buff_C9 <= data;
            8'hCA: ram_buff_CA <= data;
            8'hCB: ram_buff_CB <= data;
            8'hCC: ram_buff_CC <= data;
            8'hCD: ram_buff_CD <= data;
            8'hCE: ram_buff_CE <= data;
            8'hCF: ram_buff_CF <= data;
            8'hD0: ram_buff_D0 <= data;
            8'hD1: ram_buff_D1 <= data;
            8'hD2: ram_buff_D2 <= data;
            8'hD3: ram_buff_D3 <= data;
            8'hD4: ram_buff_D4 <= data;
            8'hD5: ram_buff_D5 <= data;
            8'hD6: ram_buff_D6 <= data;
            8'hD7: ram_buff_D7 <= data;
            8'hD8: ram_buff_D8 <= data;
            8'hD9: ram_buff_D9 <= data;
            8'hDA: ram_buff_DA <= data;
            8'hDB: ram_buff_DB <= data;
            8'hDC: ram_buff_DC <= data;
            8'hDD: ram_buff_DD <= data;
            8'hDE: ram_buff_DE <= data;
            8'hDF: ram_buff_DF <= data;
            8'hE0: ram_buff_E0 <= data;
            8'hE1: ram_buff_E1 <= data;
            8'hE2: ram_buff_E2 <= data;
            8'hE3: ram_buff_E3 <= data;
            8'hE4: ram_buff_E4 <= data;
            8'hE5: ram_buff_E5 <= data;
            8'hE6: ram_buff_E6 <= data;
            8'hE7: ram_buff_E7 <= data;
            8'hE8: ram_buff_E8 <= data;
            8'hE9: ram_buff_E9 <= data;
            8'hEA: ram_buff_EA <= data;
            8'hEB: ram_buff_EB <= data;
            8'hEC: ram_buff_EC <= data;
            8'hED: ram_buff_ED <= data;
            8'hEE: ram_buff_EE <= data;
            8'hEF: ram_buff_EF <= data;
            8'hF0: ram_buff_F0 <= data;
            8'hF1: ram_buff_F1 <= data;
            8'hF2: ram_buff_F2 <= data;
            8'hF3: ram_buff_F3 <= data;
            8'hF4: ram_buff_F4 <= data;
            8'hF5: ram_buff_F5 <= data;
            8'hF6: ram_buff_F6 <= data;
            8'hF7: ram_buff_F7 <= data;
            8'hF8: ram_buff_F8 <= data;
            8'hF9: ram_buff_F9 <= data;
            8'hFA: ram_buff_FA <= data;
            8'hFB: ram_buff_FB <= data;
            8'hFC: ram_buff_FC <= data;
            8'hFD: ram_buff_FD <= data;
            8'hFE: ram_buff_FE <= data;
            8'hFF: ram_buff_FF <= data;           
            endcase
        end
 end   
    
 always @(posedge clock)begin
         if(aclr)begin
         q <= 45'h000000000000;
         end
         else if(rden)begin
             case(rdaddress)
             8'h00: q <= ram_buff_00;
             8'h01: q <= ram_buff_01;
             8'h02: q <= ram_buff_02;
             8'h03: q <= ram_buff_03;
             8'h04: q <= ram_buff_04;
             8'h05: q <= ram_buff_05;
             8'h06: q <= ram_buff_06;
             8'h07: q <= ram_buff_07;
             8'h08: q <= ram_buff_08;
             8'h09: q <= ram_buff_09;
             8'h0A: q <= ram_buff_0A;
             8'h0B: q <= ram_buff_0B;
             8'h0C: q <= ram_buff_0C;
             8'h0D: q <= ram_buff_0D;
             8'h0E: q <= ram_buff_0E;
             8'h0F: q <= ram_buff_0F;
             8'h10: q <= ram_buff_10;
             8'h11: q <= ram_buff_11;
             8'h12: q <= ram_buff_12;
             8'h13: q <= ram_buff_13;
             8'h14: q <= ram_buff_14;
             8'h15: q <= ram_buff_15;
             8'h16: q <= ram_buff_16;
             8'h17: q <= ram_buff_17;
             8'h18: q <= ram_buff_18;
             8'h19: q <= ram_buff_19;
             8'h1A: q <= ram_buff_1A;
             8'h1B: q <= ram_buff_1B;
             8'h1C: q <= ram_buff_1C;
             8'h1D: q <= ram_buff_1D;
             8'h1E: q <= ram_buff_1E;
             8'h1F: q <= ram_buff_1F;
             8'h20: q <= ram_buff_20;
             8'h21: q <= ram_buff_21;
             8'h22: q <= ram_buff_22;
             8'h23: q <= ram_buff_23;
             8'h24: q <= ram_buff_24;
             8'h25: q <= ram_buff_25;
             8'h26: q <= ram_buff_26;
             8'h27: q <= ram_buff_27;
             8'h28: q <= ram_buff_28;
             8'h29: q <= ram_buff_29;
             8'h2A: q <= ram_buff_2A;
             8'h2B: q <= ram_buff_2B;
             8'h2C: q <= ram_buff_2C;
             8'h2D: q <= ram_buff_2D;
             8'h2E: q <= ram_buff_2E;
             8'h2F: q <= ram_buff_2F;
             8'h30: q <= ram_buff_30;
             8'h31: q <= ram_buff_31;
             8'h32: q <= ram_buff_32;
             8'h33: q <= ram_buff_33;
             8'h34: q <= ram_buff_34;
             8'h35: q <= ram_buff_35;
             8'h36: q <= ram_buff_36;
             8'h37: q <= ram_buff_37;
             8'h38: q <= ram_buff_38;
             8'h39: q <= ram_buff_39;
             8'h3A: q <= ram_buff_3A;
             8'h3B: q <= ram_buff_3B;
             8'h3C: q <= ram_buff_3C;
             8'h3D: q <= ram_buff_3D;
             8'h3E: q <= ram_buff_3E;
             8'h3F: q <= ram_buff_3F;
             8'h40: q <= ram_buff_40;
             8'h41: q <= ram_buff_41;
             8'h42: q <= ram_buff_42;
             8'h43: q <= ram_buff_43;
             8'h44: q <= ram_buff_44;
             8'h45: q <= ram_buff_45;
             8'h46: q <= ram_buff_46;
             8'h47: q <= ram_buff_47;
             8'h48: q <= ram_buff_48;
             8'h49: q <= ram_buff_49;
             8'h4A: q <= ram_buff_4A;
             8'h4B: q <= ram_buff_4B;
             8'h4C: q <= ram_buff_4C;
             8'h4D: q <= ram_buff_4D;
             8'h4E: q <= ram_buff_4E;
             8'h4F: q <= ram_buff_4F;
             8'h50: q <= ram_buff_50;
             8'h51: q <= ram_buff_51;
             8'h52: q <= ram_buff_52;
             8'h53: q <= ram_buff_53;
             8'h54: q <= ram_buff_54;
             8'h55: q <= ram_buff_55;
             8'h56: q <= ram_buff_56;
             8'h57: q <= ram_buff_57;
             8'h58: q <= ram_buff_58;
             8'h59: q <= ram_buff_59;
             8'h5A: q <= ram_buff_5A;
             8'h5B: q <= ram_buff_5B;
             8'h5C: q <= ram_buff_5C;
             8'h5D: q <= ram_buff_5D;
             8'h5E: q <= ram_buff_5E;
             8'h5F: q <= ram_buff_5F;
             8'h60: q <= ram_buff_60;
             8'h61: q <= ram_buff_61;
             8'h62: q <= ram_buff_62;
             8'h63: q <= ram_buff_63;
             8'h64: q <= ram_buff_64;
             8'h65: q <= ram_buff_65;
             8'h66: q <= ram_buff_66;
             8'h67: q <= ram_buff_67;
             8'h68: q <= ram_buff_68;
             8'h69: q <= ram_buff_69;
             8'h6A: q <= ram_buff_6A;
             8'h6B: q <= ram_buff_6B;
             8'h6C: q <= ram_buff_6C;
             8'h6D: q <= ram_buff_6D;
             8'h6E: q <= ram_buff_6E;
             8'h6F: q <= ram_buff_6F;
             8'h70: q <= ram_buff_70;
             8'h71: q <= ram_buff_71;
             8'h72: q <= ram_buff_72;
             8'h73: q <= ram_buff_73;
             8'h74: q <= ram_buff_74;
             8'h75: q <= ram_buff_75;
             8'h76: q <= ram_buff_76;
             8'h77: q <= ram_buff_77;
             8'h78: q <= ram_buff_78;
             8'h79: q <= ram_buff_79;
             8'h7A: q <= ram_buff_7A;
             8'h7B: q <= ram_buff_7B;
             8'h7C: q <= ram_buff_7C;
             8'h7D: q <= ram_buff_7D;
             8'h7E: q <= ram_buff_7E;
             8'h7F: q <= ram_buff_7F;
             8'h80: q <= ram_buff_80;
             8'h81: q <= ram_buff_81;
             8'h82: q <= ram_buff_82;
             8'h83: q <= ram_buff_83;
             8'h84: q <= ram_buff_84;
             8'h85: q <= ram_buff_85;
             8'h86: q <= ram_buff_86;
             8'h87: q <= ram_buff_87;
             8'h88: q <= ram_buff_88;
             8'h89: q <= ram_buff_89;
             8'h8A: q <= ram_buff_8A;
             8'h8B: q <= ram_buff_8B;
             8'h8C: q <= ram_buff_8C;
             8'h8D: q <= ram_buff_8D;
             8'h8E: q <= ram_buff_8E;
             8'h8F: q <= ram_buff_8F;
             8'h90: q <= ram_buff_90;
             8'h91: q <= ram_buff_91;
             8'h92: q <= ram_buff_92;
             8'h93: q <= ram_buff_93;
             8'h94: q <= ram_buff_94;
             8'h95: q <= ram_buff_95;
             8'h96: q <= ram_buff_96;
             8'h97: q <= ram_buff_97;
             8'h98: q <= ram_buff_98;
             8'h99: q <= ram_buff_99;
             8'h9A: q <= ram_buff_9A;
             8'h9B: q <= ram_buff_9B;
             8'h9C: q <= ram_buff_9C;
             8'h9D: q <= ram_buff_9D;
             8'h9E: q <= ram_buff_9E;
             8'h9F: q <= ram_buff_9F;
             8'hA0: q <= ram_buff_A0;
             8'hA1: q <= ram_buff_A1;
             8'hA2: q <= ram_buff_A2;
             8'hA3: q <= ram_buff_A3;
             8'hA4: q <= ram_buff_A4;
             8'hA5: q <= ram_buff_A5;
             8'hA6: q <= ram_buff_A6;
             8'hA7: q <= ram_buff_A7;
             8'hA8: q <= ram_buff_A8;
             8'hA9: q <= ram_buff_A9;
             8'hAA: q <= ram_buff_AA;
             8'hAB: q <= ram_buff_AB;
             8'hAC: q <= ram_buff_AC;
             8'hAD: q <= ram_buff_AD;
             8'hAE: q <= ram_buff_AE;
             8'hAF: q <= ram_buff_AF;
             8'hB0: q <= ram_buff_B0;
             8'hB1: q <= ram_buff_B1;
             8'hB2: q <= ram_buff_B2;
             8'hB3: q <= ram_buff_B3;
             8'hB4: q <= ram_buff_B4;
             8'hB5: q <= ram_buff_B5;
             8'hB6: q <= ram_buff_B6;
             8'hB7: q <= ram_buff_B7;
             8'hB8: q <= ram_buff_B8;
             8'hB9: q <= ram_buff_B9;
             8'hBA: q <= ram_buff_BA;
             8'hBB: q <= ram_buff_BB;
             8'hBC: q <= ram_buff_BC;
             8'hBD: q <= ram_buff_BD;
             8'hBE: q <= ram_buff_BE;
             8'hBF: q <= ram_buff_BF;
             8'hC0: q <= ram_buff_C0;
             8'hC1: q <= ram_buff_C1;
             8'hC2: q <= ram_buff_C2;
             8'hC3: q <= ram_buff_C3;
             8'hC4: q <= ram_buff_C4;
             8'hC5: q <= ram_buff_C5;
             8'hC6: q <= ram_buff_C6;
             8'hC7: q <= ram_buff_C7;
             8'hC8: q <= ram_buff_C8;
             8'hC9: q <= ram_buff_C9;
             8'hCA: q <= ram_buff_CA;
             8'hCB: q <= ram_buff_CB;
             8'hCC: q <= ram_buff_CC;
             8'hCD: q <= ram_buff_CD;
             8'hCE: q <= ram_buff_CE;
             8'hCF: q <= ram_buff_CF;
             8'hD0: q <= ram_buff_D0;
             8'hD1: q <= ram_buff_D1;
             8'hD2: q <= ram_buff_D2;
             8'hD3: q <= ram_buff_D3;
             8'hD4: q <= ram_buff_D4;
             8'hD5: q <= ram_buff_D5;
             8'hD6: q <= ram_buff_D6;
             8'hD7: q <= ram_buff_D7;
             8'hD8: q <= ram_buff_D8;
             8'hD9: q <= ram_buff_D9;
             8'hDA: q <= ram_buff_DA;
             8'hDB: q <= ram_buff_DB;
             8'hDC: q <= ram_buff_DC;
             8'hDD: q <= ram_buff_DD;
             8'hDE: q <= ram_buff_DE;
             8'hDF: q <= ram_buff_DF;
             8'hE0: q <= ram_buff_E0;
             8'hE1: q <= ram_buff_E1;
             8'hE2: q <= ram_buff_E2;
             8'hE3: q <= ram_buff_E3;
             8'hE4: q <= ram_buff_E4;
             8'hE5: q <= ram_buff_E5;
             8'hE6: q <= ram_buff_E6;
             8'hE7: q <= ram_buff_E7;
             8'hE8: q <= ram_buff_E8;
             8'hE9: q <= ram_buff_E9;
             8'hEA: q <= ram_buff_EA;
             8'hEB: q <= ram_buff_EB;
             8'hEC: q <= ram_buff_EC;
             8'hED: q <= ram_buff_ED;
             8'hEE: q <= ram_buff_EE;
             8'hEF: q <= ram_buff_EF;
             8'hF0: q <= ram_buff_F0;
             8'hF1: q <= ram_buff_F1;
             8'hF2: q <= ram_buff_F2;
             8'hF3: q <= ram_buff_F3;
             8'hF4: q <= ram_buff_F4;
             8'hF5: q <= ram_buff_F5;
             8'hF6: q <= ram_buff_F6;
             8'hF7: q <= ram_buff_F7;
             8'hF8: q <= ram_buff_F8;
             8'hF9: q <= ram_buff_F9;
             8'hFA: q <= ram_buff_FA;
             8'hFB: q <= ram_buff_FB;
             8'hFC: q <= ram_buff_FC;
             8'hFD: q <= ram_buff_FD;
             8'hFE: q <= ram_buff_FE;
             8'hFF: q <= ram_buff_FF;          
             endcase
         end
  end   
     
endmodule
