
`timescale 1ns / 1ps
module F_normal_t10_next_Rom4(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[159:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 160'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h13: rd_q <= 160'b1110011110000110011010010000010111111000100110111010010001001110101011001010101100110111000011010101010100010101101011100110110001111010000101111101110010000100;
			5'h12: rd_q <= 160'b1111101010000010011011111111011001111001011100011100001001110100110110000001001100101110111001110101111100010011100101101010011111100110010000010101000110011000;
			5'h11: rd_q <= 160'b1011001010011011010111100100011101111110100110000000000100001001110000000001101101101000110000100001000100110101000111010110001011110000100011111101110011010110;
			5'h10: rd_q <= 160'b0101101110100100111011100011111001110101000011010011001001001011000011001010001000001110111001111110001011000111000000110011011110110111100110001000001110111111;
			5'h0f: rd_q <= 160'b1100011010000001101011000110001011101011110111010001000010111001001001110001111101101110110100111111101011010110110101011001100000100001110111101100110111110110;
			5'h0e: rd_q <= 160'b1111000000011111100111101001011010110000011011011101111001010000100011001001010110010011001000101011010111010011101000011100111100010111101101010101000010101001;
			5'h0d: rd_q <= 160'b0101000001001001110100011110000100110001110011010001010000010011000110010110001001011101101111001001101111111101100010010011000001100000101111100001000001000011;
			5'h0c: rd_q <= 160'b1110100000110100101011010010001101100000101000101001111010000010010011010011100111011000000000101100011111010110010111011111111111001101000011110100111010100100;
			5'h0b: rd_q <= 160'b0101000101000010101101110110100010111111000111000101001001000100001001000010001000100101110010110001011001111110000101000110010000101111000010101100101100001101;
			5'h0a: rd_q <= 160'b0000000101000010000011110000110101010011101111101001010101000101101010111010010111110110000110010110011011100111111001101011110000011011010000010110101110011011;
			5'h09: rd_q <= 160'b0001111011010111000101000101101111000100010000111101100000110011010011110011110101101011011011101110100000100111011000110111101111001101100001010111100001011011;
			5'h08: rd_q <= 160'b1101001110111101001100101101001111010010011100101110101101110010000110010100011011100010100011100001101100000011110111011101111001100110111110110100000001001101;
			5'h07: rd_q <= 160'b0100010100010011100111100000011000101000101100011011111000000111011111011110110110011101111101010101111110001100101100010110101001111010100100001100111000010011;
			5'h06: rd_q <= 160'b0111000010110011111100011101001010110111011001111111100010100001011000011010101000001010010111101010100111000111111100100111111111010110110000111101110101111100;
			5'h05: rd_q <= 160'b1010011101101000100000101001001000000110010010001010001000010010010100111011100011000010110111101100000000011100001000010010000000100011111000001100111000011010;
			5'h04: rd_q <= 160'b0000001010000001111100111111011011100100000001010101101010001101110011010101000000010000101110111000010100100011001011010111000111011110111111110010001001101110;
			5'h03: rd_q <= 160'b0100001010111010010000101110000110101100100000110111011011010001000011001011110010100111101100000010101111000110010110101100001110101001001000111110110011000001;
			5'h02: rd_q <= 160'b0101100001100001000110011110110010011110110111011011001000000100111001001110110011010101011011010110011011101111010110011000100010010111011100111000110001111111;
			5'h01: rd_q <= 160'b0000101111110111110110100000011001111001100100000000111000110101010010000110100000110001011101011111010011111000100000111110001011110010010101101101101011111100;
			5'h00: rd_q <= 160'b0010111010110101000110111010010001010010010000101101111000010011000001110111101100011110101100110001001110001101010010100110111000001001111101001111001100011011;
		default:rd_q <= 160'b0;
		endcase
	end
end

endmodule
