
`timescale 1ns / 1ps
module F_normal_t8_next_Rom1(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[127:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 128'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h0f: rd_q <= 128'b01101010001100110100111110010000010101110101101100011111110011000101111011110100111100100100011101111101010100100111000000011100;
			5'h0e: rd_q <= 128'b01111011001100001111001000110000110111010100010001010001001001011100101100100110111010110100100001111101000001001101011101101001;
			5'h0d: rd_q <= 128'b11000010011111111101100011111010110000000000101110110011101111000011010100111010101100110111010110011111110100100111111100101011;
			5'h0c: rd_q <= 128'b00100000111010000011010101000100000011011011011110010100110111100101110010100000100101010001001011011101110101111110001000110101;
			5'h0b: rd_q <= 128'b11010011010011011000111011010010101011101001001101010101100011111001011100100001110110001111011010000010010110010101100100011011;
			5'h0a: rd_q <= 128'b00001111011011000111001100111110000110111010001001000100001011010101011111000101110010111100101100111111001101111100110100011010;
			5'h09: rd_q <= 128'b01001011101111101010010001000001110111110110101001001110100110101010001001001101010010111110010000000011110100000011111001011011;
			5'h08: rd_q <= 128'b01100101110001111100111110000100110111111000100010100010111110100001110000000100010101010001111101010000111001000011010001100001;
			5'h07: rd_q <= 128'b00011011010000011101100100010101110100000101010000100011001011101101110011011010111010110000110111011101111100010011000111110011;
			5'h06: rd_q <= 128'b01011101110010001111111011000011101010101100000101110000100010000000110011011110001001011101010011101000001110010110001101100011;
			5'h05: rd_q <= 128'b10010011011001000011101100100000110001111101101100011101101100000000000001011010111110010000010100010100111111001101011100001110;
			5'h04: rd_q <= 128'b11101001010110001001101110100100001010001111100001100001100110000000111001010101101100011010101011100010100011001101111001100011;
			5'h03: rd_q <= 128'b10010011110100001010101101000101101000000101100100100100101000010001000001011000011100101001000101101010111101100110001010110011;
			5'h02: rd_q <= 128'b00110111011100110010000000100001101011011110101001100010010000111101110111100110010101010000101000001001110111000001010000101100;
			5'h01: rd_q <= 128'b01010100111110001100011001110011010100101100010110101000010011010111110001100010101111000101110101010001100011011111110100000100;
			5'h00: rd_q <= 128'b10111000101000100001110010001111100011111100101001010100000000000110101110001110001110110101000110101101011100100011101011011000;
		default:rd_q <= 128'b0;
		endcase
	end
end

endmodule
