`timescale 1ns / 1ps
module F_short_t12_next_Rom7(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[167:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 168'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h14: rd_q <= 168'b010000100000001000011010101000011100000000000111111101101110010011011000010110011000011111111111011000110011011101010001100011100101001101111001000001111010011101111101;
			5'h13: rd_q <= 168'b000111111110011101011001101100100111010111010101010010010010100110001010010101011110111011101000101010110101100100010110101000010000000011011110010100000110110110001011;
			5'h12: rd_q <= 168'b111001010010101111100111000100011011011000111010010011010010001001001101100000100011000011000010001010100001011101011100001110001011001101001011010111011101110000001010;
			5'h11: rd_q <= 168'b000000100111001110101001100001010011111000011001101001011000100000001000000101011010010100100111110100001110011100001110011010100110000011010110000101000011000011000100;
			5'h10: rd_q <= 168'b101101000011101111111100111101110100110011111010001010010100110000011000011100001010011011110111001001110110010001010001010001100000000011010111010010001110000011000010;
			5'h0f: rd_q <= 168'b011100111100000011011010011100010110100101010111000111100000111100100001101001100101100001111110110110111010110010101100000100001111010100001110111011101110001100011001;
			5'h0e: rd_q <= 168'b100000101000011100110010000011101001011001000001110101010111101001010100010101101101001100010100000001101000010010101000011100010111001010011010010011111010000110111101;
			5'h0d: rd_q <= 168'b111010000101011100001000010101001100010010010111000001101110010111001001110101001100011010011010101010101101100111001110000001011110101000000011100001011100000010001110;
			5'h0c: rd_q <= 168'b111001001001011100010110011100010100011101011100110000001000111100010100111011011010001001100001110100010111000001010000011110110011101110010011001011111011111100101011;
			5'h0b: rd_q <= 168'b110011001011100010110001011111001000111111110001001110001111100101001110100111101111100111111111100011111011110011100110000110111110111100100101111001100111001001011000;
			5'h0a: rd_q <= 168'b100100101110101000011100100000011010111001010011011111010001110100110001011001001000111010101000101111010100010011001111011111100010011001010010100011101010110101010000;
			5'h09: rd_q <= 168'b000101000010011011111001000011011111110011010010101011010101010001001111111100000101110000110110001111101101010110001101011111011011110100001100101010011110011001101101;
			5'h08: rd_q <= 168'b010110011101010100100010000001010101000101100110100110101111111000100011000001111001110101101001101011011100111100011011000001000011110010110001001100110000100000001011;
			5'h07: rd_q <= 168'b010000001100110101001101111000011110101011111001000011111011101100001100001000101010011101110101000110000101011110000111101000110000111100100000111010011111100101101101;
			5'h06: rd_q <= 168'b010110011000000111001001101100011011110101110000101100010101110011001100010001000100111110010010111011101110100110011001000011101110001000000011000111110100100000010100;
			5'h05: rd_q <= 168'b000001010111010010000101000011011110111011100010010011110011101100001000011111000000101001100001101101110111010011011011111101011011111000101000101111011100010101111000;
			5'h04: rd_q <= 168'b000111101110101101101110000111001100111000101100011000110111001011000000101010011101100011101110101111001110101111011001101100000101011100000001101011100110000101100101;
			5'h03: rd_q <= 168'b110111110100110101011000101100111110111111110100000101100011110010011111011000111110110000000100101000011110111010011111011110100000111111001100011011100010110001101110;
			5'h02: rd_q <= 168'b100111110001100001100110010001101010111101111101101001110110100000100011001111011000011011011000001110100000100111010010100001001100111010001000111110110010011001000110;
			5'h01: rd_q <= 168'b100101010000001000111010111100001110010010000011010100011100110111011110111000010100010011101110101011011010011001010001000100000101000111011100110000100000011100101100;
			5'h00: rd_q <= 168'b010010011000011001010000001000101001100110001010110001010100001100101001110010111110100101101100010011111100100000011111100111010000111010001111000010010110011110010110;
		default:rd_q <= 168'b0;
		endcase
	end
end

endmodule
