
`timescale 1ns / 1ps
module F_normal_t10_next_Rom2(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[159:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 160'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h13: rd_q <= 160'b1010101111001111011010100101101011100000111101011010100100001010001100001101000010011001110000110100011011111111010000010011000001011010111111001000001000000111;
			5'h12: rd_q <= 160'b1101111111011111011100011001010011100111010111000011000111100011111000100011000011111110011010110110111011100111101000100001111000101011101001101011011001110111;
			5'h11: rd_q <= 160'b1110110011110110000011010110101111111001011100100010101111111000000000111100010111011010010100111010011111100101001001010111010100011110111111011101001101000010;
			5'h10: rd_q <= 160'b0111110111011110000000101100001011010101101111011101111011000011101100110101110000000111001100100111101010000100101001001010000110110000000000110101111011110001;
			5'h0f: rd_q <= 160'b0010111111010000011111111100011010101101111011110111101011010100000111100000000111111110101110011111100111110010101011101110000100110101110110001100011111001111;
			5'h0e: rd_q <= 160'b1111010110101000101101000001011111000011001011000100000101110010101100000010101000001001011111001100010111100111011111111011110111101100011101101011001010110011;
			5'h0d: rd_q <= 160'b0101001001101010111111011011111111000110101111010100011110100011111001000101110101001010010111111001111001101110100011001011111011101100100110010001000100000001;
			5'h0c: rd_q <= 160'b1001010100000100011110101100000010000000000100010100001000111001101101101001101100100101111111010000110111110000100011110111111010000110100111101100101010000111;
			5'h0b: rd_q <= 160'b0101011001000111011001111001100111111101111110000101111011111111000100010101110010101011100000011010100001100000111110011110111111010010010010100111110000111001;
			5'h0a: rd_q <= 160'b0000010100001000001111000011010101001110111110100101010100010110101011101001011111011000011001011001101110011111100110101111000001101101000001011010111001101100;
			5'h09: rd_q <= 160'b0111101101011100010100010110111100010001000011110110000011001101001111001111010110101101101110111010000010011101100011011110111100110110000101011110000101101100;
			5'h08: rd_q <= 160'b0111101100100010000001010000001001001011010100001001010111111000111001110110011111001111110011100111111010100110100011111111100000101001010011101111000100100011;
			5'h07: rd_q <= 160'b0000011100000011110000100010001110100011010011111110111111110010011101100110001001001011011110001000111110101010011011011101011010000100001000100110100001000001;
			5'h06: rd_q <= 160'b1101000110000010011111010111000111011100000101101111010101101010000001110111110000010101110101110101011010000111011000011000000000110101011011100010010111111101;
			5'h05: rd_q <= 160'b1011101100111001011111100011111000011010001100001010011110010110010011010100101101110010001000001110001101000001110101000111111001010011010000011001100001110010;
			5'h04: rd_q <= 160'b0000101000000111110011111101101110010000000101010110101000110111001101010100000001000010111011100001010010001100101101011100011101111011111111001000100110111000;
			5'h03: rd_q <= 160'b0001100110100100101100011011110110110011100001001100110010101011101100110010011010100010011011010101111010000001110000110111000111001010111011101110001100001001;
			5'h02: rd_q <= 160'b0111001011001001110111011000100101111010111111111101111111111100000100100110011101101001000110000110101000100101110011100101110100110011101011110110000111110001;
			5'h01: rd_q <= 160'b0010111111011111011010000001100111100110010000000011100011010101001000011010000011000101110101111101001111100010000011111000101111001001010110110110101111110000;
			5'h00: rd_q <= 160'b1011101011010100011011101001000101001001000010110111100001001100000111011110110001111010110011000100111000110101001010011011100000100111110100111100110001101100;
		default:rd_q <= 160'b0;
		endcase
	end
end

endmodule
