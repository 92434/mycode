`timescale 1ns / 1ps
module F_normal_t12_next_Rom0(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b111001111010101001000000011001101110111110100001111000101100000010010001000100001010110000111011000110110011010011110011000010100011100010001010001110100010000111000001011100000110010001110010;
			5'h16: rd_q <= 192'b100001011000100110001111000111101101011000101110000101111011110100000000011111101011011101111110100100110000110010111100111000011110001010001100011000010000010110100011001101011110110101110111;
			5'h15: rd_q <= 192'b110011100001101101001000011110111010111111110000010100100101110110010000000000011000010100101110111010111110010110101000000011111000111101000000111000001011001001010100001100010110001100010011;
			5'h14: rd_q <= 192'b111011000111001001010000101010101001101111101000110001111110011001000010011111110100000111110100110001101110111101000100001000001111100111011010101101000010111010100101101111111111000100101100;
			5'h13: rd_q <= 192'b100000010010000110101100000011001011011010011001110101100000010100100000011000010001111101000010011010000110010000010011000000101011000101101011010010001011001000100101010111110110000001010000;
			5'h12: rd_q <= 192'b000111000111010001101001101000001101000101000010101001011000111000010111000000100111010010011000001000010000111011111010011100100100010110100000001011000000110010001010000010110101001111101110;
			5'h11: rd_q <= 192'b010100100111010101110111010011010001110111011110011111111011000011110110001101011010110100110001100001001010010110100001100010001101111000010101000011011100100100101101010011100110111001001010;
			5'h10: rd_q <= 192'b111001000110011010011100000100000011100100000010101110110011010000100011101000101101101100100110110001101101110010000101011001111001100010110110000001111100010010001111010110001110101110001101;
			5'h0f: rd_q <= 192'b011111001000010010110110001010011100010011001100101011100011001011110100100110001101111101011101011011001101100110000011110101101100110000100100000111001100000101111011101000101000110001011101;
			5'h0e: rd_q <= 192'b100001110100001101011100011010011100111101100100101111101011111101110001011111010101110011100101011011110010000111101011101110110000001011101011111100111011111110000111000010000001111011000110;
			5'h0d: rd_q <= 192'b010111001001010011100100011111101011101000111010010001111000011111001110010000101101100011011010010010000101100011000001101010011011010011011010111001011011010010000010010101000110101101000000;
			5'h0c: rd_q <= 192'b011100111000100110110100110101110000100101101010110010110010011111001111010001100001010011000101010101111101001000100001010001001011010111110001110001111111010101010100001110100110011001010010;
			5'h0b: rd_q <= 192'b010110110101110101111100100101010011001110000001010001101110010001010010011101000110011011110011101100001011100110010101111110110001101010101001101011100101000111000110100011001101101000011011;
			5'h0a: rd_q <= 192'b001111001101110101100010111001110100111111000111001100101010111001000111111110001011100111100001011101111111111010011000111001010001100001101111010010100110101111101011000101100011011110111100;
			5'h09: rd_q <= 192'b000010010111101100101011011001111011111011001000110101100000100010100011110111100111011100011011100010000001110100010110001100000001011101010100100111010011100101111001111101111001001101010011;
			5'h08: rd_q <= 192'b100111110110000000010000111110101111000000101001000011100000001001011111110001001100100000011011011111100001011011000101000110111101101000000111101111010100001111001110001010100000010111100101;
			5'h07: rd_q <= 192'b000000010101000000110100100100000011011100101111011010101100101110000011011111011110010110010000011011010100100001111111001000110000111110101011000100111100100100000000010011001100101011001101;
			5'h06: rd_q <= 192'b000011111011010010100000101100100011001100010010011100101000001101000011101100000101011001111110010101111110100001101110101010011001010011110110000111001100010110010110100101011010101001000101;
			5'h05: rd_q <= 192'b001110000010101001110000001110011100010000000100001010010000011100100110001001011011101000000000110011101010110010111101010010100011001111000111011011001110000011110110010010000110110001111110;
			5'h04: rd_q <= 192'b110110101101101100000001000011011100000101001110000101101100010010110100101111100110010101011110111010011000001000010111001000011000010110111101000010101111110011011000110101000111011110110000;
			5'h03: rd_q <= 192'b010101100001000000100011001001110001110000001101111110111001111010111010010110101101011011110001011101101101100001011001001100011111010011110011011010011101011001010100000100101111001111011100;
			5'h02: rd_q <= 192'b101001001000010000010110011010100101110100000010011101111101000101101110111111110000010001011100110010000111111110000110101111000110100101010101101010001010001110010101110111001101100011000000;
			5'h01: rd_q <= 192'b100101001101101111100100010000111111001000101100000100011101011100001000111101100000010100100010110010100110011011110101000010011001100010100110011100101001100110000010010111011000101010010011;
			5'h00: rd_q <= 192'b000010111000001011010000011000000100110000010100111110010110010101011001111101110001101001001111110100011111101000110100011101111100011101000111011010001001110101001111000110011111100110110111;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
