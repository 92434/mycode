`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2015/08/30 16:10:39
// Design Name: 
// Module Name: total_yu_Q_360_rom_txt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module total_yu_Q_360_rom_txt(
    input [12:0] address,
    input clock,
    input rden,
    output reg [7:0] q
    );
    
    always @(posedge clock)begin
        if(rden == 1'b1)begin
            case(address)
            12'h0000:q <= 8'h74;
            12'h0001:q <= 8'h35;
            12'h0002:q <= 8'h3C;
            12'h0003:q <= 8'h68;
            12'h0004:q <= 8'h3A;
            12'h0005:q <= 8'h0F;
            12'h0006:q <= 8'h10;
            12'h0007:q <= 8'h00;
            12'h0008:q <= 8'h1D;
            12'h0009:q <= 8'h59;
            12'h000A:q <= 8'h2A;
            12'h000B:q <= 8'h6C;
            12'h000C:q <= 8'hFF;
            12'h000D:q <= 8'h54;
            12'h000E:q <= 8'h58;
            12'h000F:q <= 8'h04;
            12'h0010:q <= 8'h67;
            12'h0011:q <= 8'h85;
            12'h0012:q <= 8'h16;
            12'h0013:q <= 8'h3E;
            12'h0014:q <= 8'h76;
            12'h0015:q <= 8'h5B;
            12'h0016:q <= 8'h75;
            12'h0017:q <= 8'h22;
            12'h0018:q <= 8'h25;
            12'h0019:q <= 8'hFF;
            12'h001A:q <= 8'h77;
            12'h001B:q <= 8'h86;
            12'h001C:q <= 8'h4A;
            12'h001D:q <= 8'h1D;
            12'h001E:q <= 8'h63;
            12'h001F:q <= 8'h2C;
            12'h0020:q <= 8'h0B;
            12'h0021:q <= 8'h47;
            12'h0022:q <= 8'h3B;
            12'h0023:q <= 8'h58;
            12'h0024:q <= 8'h0F;
            12'h0025:q <= 8'h37;
            12'h0026:q <= 8'hFF;
            12'h0027:q <= 8'h72;
            12'h0028:q <= 8'h40;
            12'h0029:q <= 8'h64;
            12'h002A:q <= 8'h7A;
            12'h002B:q <= 8'h3B;
            12'h002C:q <= 8'h83;
            12'h002D:q <= 8'h26;
            12'h002E:q <= 8'h84;
            12'h002F:q <= 8'h1B;
            12'h0030:q <= 8'h53;
            12'h0031:q <= 8'h72;
            12'h0032:q <= 8'h5E;
            12'h0033:q <= 8'hFF;
            12'h0034:q <= 8'h48;
            12'h0035:q <= 8'h24;
            12'h0036:q <= 8'h32;
            12'h0037:q <= 8'h56;
            12'h0038:q <= 8'h34;
            12'h0039:q <= 8'h1B;
            12'h003A:q <= 8'h4A;
            12'h003B:q <= 8'h7E;
            12'h003C:q <= 8'h6D;
            12'h003D:q <= 8'h05;
            12'h003E:q <= 8'h50;
            12'h003F:q <= 8'h1F;
            12'h0040:q <= 8'hFF;
            12'h0041:q <= 8'h28;
            12'h0042:q <= 8'h53;
            12'h0043:q <= 8'h06;
            12'h0044:q <= 8'h19;
            12'h0045:q <= 8'h1F;
            12'h0046:q <= 8'h2D;
            12'h0047:q <= 8'h68;
            12'h0048:q <= 8'h06;
            12'h0049:q <= 8'h4D;
            12'h004A:q <= 8'h83;
            12'h004B:q <= 8'h49;
            12'h004C:q <= 8'h80;
            12'h004D:q <= 8'hFF;
            12'h004E:q <= 8'h71;
            12'h004F:q <= 8'h6C;
            12'h0050:q <= 8'h2E;
            12'h0051:q <= 8'h18;
            12'h0052:q <= 8'h50;
            12'h0053:q <= 8'h1E;
            12'h0054:q <= 8'h6F;
            12'h0055:q <= 8'h02;
            12'h0056:q <= 8'h24;
            12'h0057:q <= 8'h41;
            12'h0058:q <= 8'h39;
            12'h0059:q <= 8'h30;
            12'h005A:q <= 8'hFF;
            12'h005B:q <= 8'h49;
            12'h005C:q <= 8'h10;
            12'h005D:q <= 8'h65;
            12'h005E:q <= 8'h82;
            12'h005F:q <= 8'h33;
            12'h0060:q <= 8'h7C;
            12'h0061:q <= 8'h2F;
            12'h0062:q <= 8'h85;
            12'h0063:q <= 8'h57;
            12'h0064:q <= 8'h1C;
            12'h0065:q <= 8'h62;
            12'h0066:q <= 8'h3C;
            12'h0067:q <= 8'hFF;
            12'h0068:q <= 8'h5A;
            12'h0069:q <= 8'h22;
            12'h006A:q <= 8'h46;
            12'h006B:q <= 8'h11;
            12'h006C:q <= 8'h55;
            12'h006D:q <= 8'h43;
            12'h006E:q <= 8'h2D;
            12'h006F:q <= 8'h18;
            12'h0070:q <= 8'h0C;
            12'h0071:q <= 8'h56;
            12'h0072:q <= 8'h13;
            12'h0073:q <= 8'h34;
            12'h0074:q <= 8'hFF;
            12'h0075:q <= 8'h84;
            12'h0076:q <= 8'h45;
            12'h0077:q <= 8'h4B;
            12'h0078:q <= 8'h12;
            12'h0079:q <= 8'h25;
            12'h007A:q <= 8'h39;
            12'h007B:q <= 8'h73;
            12'h007C:q <= 8'h71;
            12'h007D:q <= 8'h2C;
            12'h007E:q <= 8'h0A;
            12'h007F:q <= 8'h27;
            12'h0080:q <= 8'h63;
            12'h0081:q <= 8'hFF;
            12'h0082:q <= 8'h0A;
            12'h0083:q <= 8'h6F;
            12'h0084:q <= 8'h07;
            12'h0085:q <= 8'h23;
            12'h0086:q <= 8'h17;
            12'h0087:q <= 8'h76;
            12'h0088:q <= 8'h79;
            12'h0089:q <= 8'h6A;
            12'h008A:q <= 8'h67;
            12'h008B:q <= 8'h64;
            12'h008C:q <= 8'h6B;
            12'h008D:q <= 8'h4B;
            12'h008E:q <= 8'hFF;
            12'h008F:q <= 8'h4F;
            12'h0090:q <= 8'h30;
            12'h0091:q <= 8'h41;
            12'h0092:q <= 8'h3D;
            12'h0093:q <= 8'h44;
            12'h0094:q <= 8'h14;
            12'h0095:q <= 8'h0E;
            12'h0096:q <= 8'h51;
            12'h0097:q <= 8'h04;
            12'h0098:q <= 8'h36;
            12'h0099:q <= 8'h21;
            12'h009A:q <= 8'h31;
            12'h009B:q <= 8'hFF;
            12'h009C:q <= 8'h59;
            12'h009D:q <= 8'h0B;
            12'h009E:q <= 8'h4D;
            12'h009F:q <= 8'h4C;
            12'h00A0:q <= 8'h5E;
            12'h00A1:q <= 8'h13;
            12'h00A2:q <= 8'h5A;
            12'h00A3:q <= 8'h43;
            12'h00A4:q <= 8'h11;
            12'h00A5:q <= 8'h2E;
            12'h00A6:q <= 8'h60;
            12'h00A7:q <= 8'h07;
            12'h00A8:q <= 8'hFF;
            12'h00A9:q <= 8'h75;
            12'h00AA:q <= 8'h42;
            12'h00AB:q <= 8'h31;
            12'h00AC:q <= 8'h80;
            12'h00AD:q <= 8'h29;
            12'h00AE:q <= 8'h66;
            12'h00AF:q <= 8'h40;
            12'h00B0:q <= 8'h33;
            12'h00B1:q <= 8'h19;
            12'h00B2:q <= 8'h03;
            12'h00B3:q <= 8'h35;
            12'h00B4:q <= 8'h29;
            12'h00B5:q <= 8'hFF;
            12'h00B6:q <= 8'h3F;
            12'h00B7:q <= 8'h0D;
            12'h00B8:q <= 8'h6B;
            12'h00B9:q <= 8'h1C;
            12'h00BA:q <= 8'h6E;
            12'h00BB:q <= 8'h02;
            12'h00BC:q <= 8'h7D;
            12'h00BD:q <= 8'h81;
            12'h00BE:q <= 8'h77;
            12'h00BF:q <= 8'h61;
            12'h00C0:q <= 8'h15;
            12'h00C1:q <= 8'h4E;
            12'h00C2:q <= 8'hFF;
            12'h00C3:q <= 8'h0C;
            12'h00C4:q <= 8'h60;
            12'h00C5:q <= 8'h3E;
            12'h00C6:q <= 8'hFF;
            12'h00C7:q <= 8'h2A;
            12'h00C8:q <= 8'h7B;
            12'h00C9:q <= 8'h7F;
            12'h00CA:q <= 8'hFF;
            12'h00CB:q <= 8'h1A;
            12'h00CC:q <= 8'h09;
            12'h00CD:q <= 8'h51;
            12'h00CE:q <= 8'hFF;
            12'h00CF:q <= 8'h52;
            12'h00D0:q <= 8'h5F;
            12'h00D1:q <= 8'h5D;
            12'h00D2:q <= 8'hFF;
            12'h00D3:q <= 8'h62;
            12'h00D4:q <= 8'h2F;
            12'h00D5:q <= 8'h27;
            12'h00D6:q <= 8'hFF;
            12'h00D7:q <= 8'h7E;
            12'h00D8:q <= 8'h73;
            12'h00D9:q <= 8'h03;
            12'h00DA:q <= 8'hFF;
            12'h00DB:q <= 8'h2B;
            12'h00DC:q <= 8'h61;
            12'h00DD:q <= 8'h78;
            12'h00DE:q <= 8'hFF;
            12'h00DF:q <= 8'h7D;
            12'h00E0:q <= 8'h38;
            12'h00E1:q <= 8'h37;
            12'h00E2:q <= 8'hFF;
            12'h00E3:q <= 8'h36;
            12'h00E4:q <= 8'h70;
            12'h00E5:q <= 8'h15;
            12'h00E6:q <= 8'hFF;
            12'h00E7:q <= 8'h08;
            12'h00E8:q <= 8'h57;
            12'h00E9:q <= 8'h20;
            12'h00EA:q <= 8'hFF;
            12'h00EB:q <= 8'h21;
            12'h00EC:q <= 8'h05;
            12'h00ED:q <= 8'h81;
            12'h00EE:q <= 8'hFF;
            12'h00EF:q <= 8'h47;
            12'h00F0:q <= 8'h79;
            12'h00F1:q <= 8'h4E;
            12'h00F2:q <= 8'hFF;
            12'h00F3:q <= 8'h69;
            12'h00F4:q <= 8'h00;
            12'h00F5:q <= 8'h26;
            12'h00F6:q <= 8'hFF;
            12'h00F7:q <= 8'h01;
            12'h00F8:q <= 8'h6D;
            12'h00F9:q <= 8'h5B;
            12'h00FA:q <= 8'hFF;
            12'h00FB:q <= 8'h0E;
            12'h00FC:q <= 8'h5C;
            12'h00FD:q <= 8'h6A;
            12'h00FE:q <= 8'hFF;
            12'h00FF:q <= 8'h1E;
            12'h0100:q <= 8'h7F;
            12'h0101:q <= 8'h14;
            12'h0102:q <= 8'hFF;
            12'h0103:q <= 8'h65;
            12'h0104:q <= 8'h54;
            12'h0105:q <= 8'h32;
            12'h0106:q <= 8'hFF;
            12'h0107:q <= 8'h74;
            12'h0108:q <= 8'h52;
            12'h0109:q <= 8'h55;
            12'h010A:q <= 8'hFF;
            12'h010B:q <= 8'h82;
            12'h010C:q <= 8'h42;
            12'h010D:q <= 8'h28;
            12'h010E:q <= 8'hFF;
            12'h010F:q <= 8'h48;
            12'h0110:q <= 8'h7A;
            12'h0111:q <= 8'h1A;
            12'h0112:q <= 8'hFF;
            12'h0113:q <= 8'h08;
            12'h0114:q <= 8'h16;
            12'h0115:q <= 8'h45;
            12'h0116:q <= 8'hFF;
            12'h0117:q <= 8'h17;
            12'h0118:q <= 8'h86;
            12'h0119:q <= 8'h20;
            12'h011A:q <= 8'hFF;
            12'h011B:q <= 8'h2B;
            12'h011C:q <= 8'h38;
            12'h011D:q <= 8'h5C;
            12'h011E:q <= 8'hFF;
            12'h011F:q <= 8'h44;
            12'h0120:q <= 8'h3A;
            12'h0121:q <= 8'h46;
            12'h0122:q <= 8'hFF;
            12'h0123:q <= 8'h4F;
            12'h0124:q <= 8'h4C;
            12'h0125:q <= 8'h3D;
            12'h0126:q <= 8'hFF;
            12'h0127:q <= 8'h12;
            12'h0128:q <= 8'h69;
            12'h0129:q <= 8'h23;
            12'h012A:q <= 8'hFF;
            12'h012B:q <= 8'h3F;
            12'h012C:q <= 8'h5F;
            12'h012D:q <= 8'h09;
            12'h012E:q <= 8'hFF;
            12'h012F:q <= 8'h5D;
            12'h0130:q <= 8'h7C;
            12'h0131:q <= 8'h0D;
            12'h0132:q <= 8'hFF;
            12'h0133:q <= 8'h7B;
            12'h0134:q <= 8'h70;
            12'h0135:q <= 8'h78;
            12'h0136:q <= 8'hFF;
            12'h0137:q <= 8'h6E;
            12'h0138:q <= 8'h66;
            12'h0139:q <= 8'h01;
            12'h013A:q <= 8'hFF;
            12'h013B:q <= 8'h1F;
            12'h013C:q <= 8'h0E;
            12'h013D:q <= 8'h10;
            12'h013E:q <= 8'h1B;
            12'h013F:q <= 8'h0F;
            12'h0140:q <= 8'h04;
            12'h0141:q <= 8'h04;
            12'h0142:q <= 8'h00;
            12'h0143:q <= 8'h07;
            12'h0144:q <= 8'h17;
            12'h0145:q <= 8'h0B;
            12'h0146:q <= 8'h1D;
            12'h0147:q <= 8'hFF;
            12'h0148:q <= 8'h23;
            12'h0149:q <= 8'h14;
            12'h014A:q <= 8'h07;
            12'h014B:q <= 8'h1A;
            12'h014C:q <= 8'h0B;
            12'h014D:q <= 8'h02;
            12'h014E:q <= 8'h13;
            12'h014F:q <= 8'h11;
            12'h0150:q <= 8'h18;
            12'h0151:q <= 8'h05;
            12'h0152:q <= 8'h10;
            12'h0153:q <= 8'h02;
            12'h0154:q <= 8'hFF;
            12'h0155:q <= 8'h0A;
            12'h0156:q <= 8'h0D;
            12'h0157:q <= 8'h18;
            12'h0158:q <= 8'h11;
            12'h0159:q <= 8'h08;
            12'h015A:q <= 8'h15;
            12'h015B:q <= 8'h22;
            12'h015C:q <= 8'h1F;
            12'h015D:q <= 8'h03;
            12'h015E:q <= 8'h19;
            12'h015F:q <= 8'h0A;
            12'h0160:q <= 8'h08;
            12'h0161:q <= 8'hFF;
            12'h0162:q <= 8'h19;
            12'h0163:q <= 8'h00;
            12'h0164:q <= 8'h05;
            12'h0165:q <= 8'h06;
            12'h0166:q <= 8'h0C;
            12'h0167:q <= 8'h1E;
            12'h0168:q <= 8'h01;
            12'h0169:q <= 8'h16;
            12'h016A:q <= 8'h23;
            12'h016B:q <= 8'h15;
            12'h016C:q <= 8'h21;
            12'h016D:q <= 8'h20;
            12'h016E:q <= 8'hFF;
            12'h016F:q <= 8'h20;
            12'h0170:q <= 8'h13;
            12'h0171:q <= 8'h09;
            12'h0172:q <= 8'hFF;
            12'h0173:q <= 8'h01;
            12'h0174:q <= 8'h12;
            12'h0175:q <= 8'h17;
            12'h0176:q <= 8'hFF;
            12'h0177:q <= 8'h1C;
            12'h0178:q <= 8'h16;
            12'h0179:q <= 8'h22;
            12'h017A:q <= 8'hFF;
            12'h017B:q <= 8'h21;
            12'h017C:q <= 8'h1D;
            12'h017D:q <= 8'h03;
            12'h017E:q <= 8'hFF;
            12'h017F:q <= 8'h0C;
            12'h0180:q <= 8'h12;
            12'h0181:q <= 8'h09;
            12'h0182:q <= 8'hFF;
            12'h0183:q <= 8'h67;
            12'h0184:q <= 8'h2F;
            12'h0185:q <= 8'h35;
            12'h0186:q <= 8'h5C;
            12'h0187:q <= 8'h33;
            12'h0188:q <= 8'h0D;
            12'h0189:q <= 8'h0E;
            12'h018A:q <= 8'h00;
            12'h018B:q <= 8'h1A;
            12'h018C:q <= 8'h4F;
            12'h018D:q <= 8'h26;
            12'h018E:q <= 8'h00;
            12'h018F:q <= 8'hFF;
            12'h0190:q <= 8'h74;
            12'h0191:q <= 8'h4A;
            12'h0192:q <= 8'h4E;
            12'h0193:q <= 8'h03;
            12'h0194:q <= 8'h5D;
            12'h0195:q <= 8'h76;
            12'h0196:q <= 8'h16;
            12'h0197:q <= 8'h38;
            12'h0198:q <= 8'h69;
            12'h0199:q <= 8'h51;
            12'h019A:q <= 8'h68;
            12'h019B:q <= 8'h1E;
            12'h019C:q <= 8'hFF;
            12'h019D:q <= 8'h31;
            12'h019E:q <= 8'h69;
            12'h019F:q <= 8'h77;
            12'h01A0:q <= 8'h40;
            12'h01A1:q <= 8'h1B;
            12'h01A2:q <= 8'h59;
            12'h01A3:q <= 8'h29;
            12'h01A4:q <= 8'h0A;
            12'h01A5:q <= 8'h3E;
            12'h01A6:q <= 8'h34;
            12'h01A7:q <= 8'h4E;
            12'h01A8:q <= 8'h0E;
            12'h01A9:q <= 8'hFF;
            12'h01AA:q <= 8'h4B;
            12'h01AB:q <= 8'h64;
            12'h01AC:q <= 8'h38;
            12'h01AD:q <= 8'h59;
            12'h01AE:q <= 8'h6D;
            12'h01AF:q <= 8'h39;
            12'h01B0:q <= 8'h75;
            12'h01B1:q <= 8'h22;
            12'h01B2:q <= 8'h75;
            12'h01B3:q <= 8'h17;
            12'h01B4:q <= 8'h49;
            12'h01B5:q <= 8'h64;
            12'h01B6:q <= 8'hFF;
            12'h01B7:q <= 8'h48;
            12'h01B8:q <= 8'h3F;
            12'h01B9:q <= 8'h1F;
            12'h01BA:q <= 8'h2B;
            12'h01BB:q <= 8'h50;
            12'h01BC:q <= 8'h35;
            12'h01BD:q <= 8'h1C;
            12'h01BE:q <= 8'h43;
            12'h01BF:q <= 8'h70;
            12'h01C0:q <= 8'h60;
            12'h01C1:q <= 8'h05;
            12'h01C2:q <= 8'h46;
            12'h01C3:q <= 8'hFF;
            12'h01C4:q <= 8'h15;
            12'h01C5:q <= 8'h23;
            12'h01C6:q <= 8'h4C;
            12'h01C7:q <= 8'h06;
            12'h01C8:q <= 8'h1A;
            12'h01C9:q <= 8'h20;
            12'h01CA:q <= 8'h2D;
            12'h01CB:q <= 8'h5F;
            12'h01CC:q <= 8'h06;
            12'h01CD:q <= 8'h42;
            12'h01CE:q <= 8'h74;
            12'h01CF:q <= 8'h3F;
            12'h01D0:q <= 8'hFF;
            12'h01D1:q <= 8'h55;
            12'h01D2:q <= 8'h66;
            12'h01D3:q <= 8'h60;
            12'h01D4:q <= 8'h26;
            12'h01D5:q <= 8'h19;
            12'h01D6:q <= 8'h4A;
            12'h01D7:q <= 8'h1E;
            12'h01D8:q <= 8'h64;
            12'h01D9:q <= 8'h02;
            12'h01DA:q <= 8'h20;
            12'h01DB:q <= 8'h39;
            12'h01DC:q <= 8'h62;
            12'h01DD:q <= 8'hFF;
            12'h01DE:q <= 8'h12;
            12'h01DF:q <= 8'h16;
            12'h01E0:q <= 8'h3D;
            12'h01E1:q <= 8'h0F;
            12'h01E2:q <= 8'h5B;
            12'h01E3:q <= 8'h74;
            12'h01E4:q <= 8'h31;
            12'h01E5:q <= 8'h6E;
            12'h01E6:q <= 8'h2A;
            12'h01E7:q <= 8'h76;
            12'h01E8:q <= 8'h4C;
            12'h01E9:q <= 8'h1B;
            12'h01EA:q <= 8'hFF;
            12'h01EB:q <= 8'h68;
            12'h01EC:q <= 8'h1A;
            12'h01ED:q <= 8'h76;
            12'h01EE:q <= 8'h3C;
            12'h01EF:q <= 8'h44;
            12'h01F0:q <= 8'h12;
            12'h01F1:q <= 8'h25;
            12'h01F2:q <= 8'h37;
            12'h01F3:q <= 8'h63;
            12'h01F4:q <= 8'h5F;
            12'h01F5:q <= 8'h25;
            12'h01F6:q <= 8'h0B;
            12'h01F7:q <= 8'hFF;
            12'h01F8:q <= 8'h09;
            12'h01F9:q <= 8'h56;
            12'h01FA:q <= 8'h0B;
            12'h01FB:q <= 8'h62;
            12'h01FC:q <= 8'h07;
            12'h01FD:q <= 8'h26;
            12'h01FE:q <= 8'h18;
            12'h01FF:q <= 8'h69;
            12'h0200:q <= 8'h6B;
            12'h0201:q <= 8'h5B;
            12'h0202:q <= 8'h59;
            12'h0203:q <= 8'h56;
            12'h0204:q <= 8'hFF;
            12'h0205:q <= 8'h14;
            12'h0206:q <= 8'h5E;
            12'h0207:q <= 8'h43;
            12'h0208:q <= 8'h28;
            12'h0209:q <= 8'h3F;
            12'h020A:q <= 8'h3A;
            12'h020B:q <= 8'h41;
            12'h020C:q <= 8'h13;
            12'h020D:q <= 8'h0D;
            12'h020E:q <= 8'h45;
            12'h020F:q <= 8'h04;
            12'h0210:q <= 8'h2E;
            12'h0211:q <= 8'hFF;
            12'h0212:q <= 8'h39;
            12'h0213:q <= 8'h2D;
            12'h0214:q <= 8'h44;
            12'h0215:q <= 8'h0D;
            12'h0216:q <= 8'h46;
            12'h0217:q <= 8'h42;
            12'h0218:q <= 8'h53;
            12'h0219:q <= 8'h15;
            12'h021A:q <= 8'h4A;
            12'h021B:q <= 8'h37;
            12'h021C:q <= 8'h0F;
            12'h021D:q <= 8'h27;
            12'h021E:q <= 8'hFF;
            12'h021F:q <= 8'h57;
            12'h0220:q <= 8'h6B;
            12'h0221:q <= 8'h6A;
            12'h0222:q <= 8'h37;
            12'h0223:q <= 8'h30;
            12'h0224:q <= 8'h73;
            12'h0225:q <= 8'h28;
            12'h0226:q <= 8'h57;
            12'h0227:q <= 8'h32;
            12'h0228:q <= 8'h2B;
            12'h0229:q <= 8'h16;
            12'h022A:q <= 8'h03;
            12'h022B:q <= 8'hFF;
            12'h022C:q <= 8'h53;
            12'h022D:q <= 8'h1D;
            12'h022E:q <= 8'h33;
            12'h022F:q <= 8'h11;
            12'h0230:q <= 8'h60;
            12'h0231:q <= 8'h1F;
            12'h0232:q <= 8'h63;
            12'h0233:q <= 8'h04;
            12'h0234:q <= 8'h6D;
            12'h0235:q <= 8'h72;
            12'h0236:q <= 8'h61;
            12'h0237:q <= 8'h53;
            12'h0238:q <= 8'hFF;
            12'h0239:q <= 8'h49;
            12'h023A:q <= 8'h46;
            12'h023B:q <= 8'h50;
            12'h023C:q <= 8'h27;
            12'h023D:q <= 8'h2B;
            12'h023E:q <= 8'h14;
            12'h023F:q <= 8'h77;
            12'h0240:q <= 8'h27;
            12'h0241:q <= 8'h6F;
            12'h0242:q <= 8'h5C;
            12'h0243:q <= 8'h0C;
            12'h0244:q <= 8'h5A;
            12'h0245:q <= 8'hFF;
            12'h0246:q <= 8'h42;
            12'h0247:q <= 8'h34;
            12'h0248:q <= 8'h2E;
            12'h0249:q <= 8'h6E;
            12'h024A:q <= 8'h23;
            12'h024B:q <= 8'h3C;
            12'h024C:q <= 8'h06;
            12'h024D:q <= 8'h45;
            12'h024E:q <= 8'h19;
            12'h024F:q <= 8'h3D;
            12'h0250:q <= 8'h3C;
            12'h0251:q <= 8'h23;
            12'h0252:q <= 8'hFF;
            12'h0253:q <= 8'h29;
            12'h0254:q <= 8'h0C;
            12'h0255:q <= 8'h71;
            12'h0256:q <= 8'h1E;
            12'h0257:q <= 8'h5E;
            12'h0258:q <= 8'h02;
            12'h0259:q <= 8'h32;
            12'h025A:q <= 8'h0B;
            12'h025B:q <= 8'h15;
            12'h025C:q <= 8'h33;
            12'h025D:q <= 8'h09;
            12'h025E:q <= 8'h67;
            12'h025F:q <= 8'hFF;
            12'h0260:q <= 8'h10;
            12'h0261:q <= 8'h3E;
            12'h0262:q <= 8'h6D;
            12'h0263:q <= 8'h17;
            12'h0264:q <= 8'h2F;
            12'h0265:q <= 8'h6F;
            12'h0266:q <= 8'h4B;
            12'h0267:q <= 8'h05;
            12'h0268:q <= 8'h1C;
            12'h0269:q <= 8'h3A;
            12'h026A:q <= 8'h47;
            12'h026B:q <= 8'h55;
            12'h026C:q <= 8'hFF;
            12'h026D:q <= 8'h05;
            12'h026E:q <= 8'h2A;
            12'h026F:q <= 8'h19;
            12'h0270:q <= 8'h32;
            12'h0271:q <= 8'h24;
            12'h0272:q <= 8'h54;
            12'h0273:q <= 8'h47;
            12'h0274:q <= 8'h49;
            12'h0275:q <= 8'h30;
            12'h0276:q <= 8'h28;
            12'h0277:q <= 8'h07;
            12'h0278:q <= 8'h2C;
            12'h0279:q <= 8'hFF;
            12'h027A:q <= 8'h4F;
            12'h027B:q <= 8'h20;
            12'h027C:q <= 8'h70;
            12'h027D:q <= 8'h0A;
            12'h027E:q <= 8'h70;
            12'h027F:q <= 8'h56;
            12'h0280:q <= 8'h58;
            12'h0281:q <= 8'h6A;
            12'h0282:q <= 8'h43;
            12'h0283:q <= 8'h57;
            12'h0284:q <= 8'h35;
            12'h0285:q <= 8'h58;
            12'h0286:q <= 8'hFF;
            12'h0287:q <= 8'h6C;
            12'h0288:q <= 8'h1D;
            12'h0289:q <= 8'h3B;
            12'h028A:q <= 8'hFF;
            12'h028B:q <= 8'h08;
            12'h028C:q <= 8'h72;
            12'h028D:q <= 8'h71;
            12'h028E:q <= 8'hFF;
            12'h028F:q <= 8'h0E;
            12'h0290:q <= 8'h08;
            12'h0291:q <= 8'h13;
            12'h0292:q <= 8'hFF;
            12'h0293:q <= 8'h04;
            12'h0294:q <= 8'h09;
            12'h0295:q <= 8'h41;
            12'h0296:q <= 8'hFF;
            12'h0297:q <= 8'h45;
            12'h0298:q <= 8'h52;
            12'h0299:q <= 8'h22;
            12'h029A:q <= 8'hFF;
            12'h029B:q <= 8'h25;
            12'h029C:q <= 8'h3B;
            12'h029D:q <= 8'h5E;
            12'h029E:q <= 8'hFF;
            12'h029F:q <= 8'h5D;
            12'h02A0:q <= 8'h4E;
            12'h02A1:q <= 8'h48;
            12'h02A2:q <= 8'hFF;
            12'h02A3:q <= 8'h02;
            12'h02A4:q <= 8'h34;
            12'h02A5:q <= 8'h50;
            12'h02A6:q <= 8'hFF;
            12'h02A7:q <= 8'h5A;
            12'h02A8:q <= 8'h3D;
            12'h02A9:q <= 8'h65;
            12'h02AA:q <= 8'hFF;
            12'h02AB:q <= 8'h41;
            12'h02AC:q <= 8'h17;
            12'h02AD:q <= 8'h36;
            12'h02AE:q <= 8'hFF;
            12'h02AF:q <= 8'h73;
            12'h02B0:q <= 8'h2C;
            12'h02B1:q <= 8'h5D;
            12'h02B2:q <= 8'hFF;
            12'h02B3:q <= 8'h5F;
            12'h02B4:q <= 8'h71;
            12'h02B5:q <= 8'h52;
            12'h02B6:q <= 8'hFF;
            12'h02B7:q <= 8'h47;
            12'h02B8:q <= 8'h65;
            12'h02B9:q <= 8'h14;
            12'h02BA:q <= 8'hFF;
            12'h02BB:q <= 8'h63;
            12'h02BC:q <= 8'h48;
            12'h02BD:q <= 8'h21;
            12'h02BE:q <= 8'hFF;
            12'h02BF:q <= 8'h6F;
            12'h02C0:q <= 8'h11;
            12'h02C1:q <= 8'h08;
            12'h02C2:q <= 8'hFF;
            12'h02C3:q <= 8'h54;
            12'h02C4:q <= 8'h01;
            12'h02C5:q <= 8'h11;
            12'h02C6:q <= 8'hFF;
            12'h02C7:q <= 8'h3B;
            12'h02C8:q <= 8'h5C;
            12'h02C9:q <= 8'h77;
            12'h02CA:q <= 8'hFF;
            12'h02CB:q <= 8'h36;
            12'h02CC:q <= 8'h4D;
            12'h02CD:q <= 8'h18;
            12'h02CE:q <= 8'hFF;
            12'h02CF:q <= 8'h52;
            12'h02D0:q <= 8'h4C;
            12'h02D1:q <= 8'h4D;
            12'h02D2:q <= 8'hFF;
            12'h02D3:q <= 8'h61;
            12'h02D4:q <= 8'h2E;
            12'h02D5:q <= 8'h40;
            12'h02D6:q <= 8'hFF;
            12'h02D7:q <= 8'h72;
            12'h02D8:q <= 8'h67;
            12'h02D9:q <= 8'h24;
            12'h02DA:q <= 8'hFF;
            12'h02DB:q <= 8'h5B;
            12'h02DC:q <= 8'h5A;
            12'h02DD:q <= 8'h1D;
            12'h02DE:q <= 8'hFF;
            12'h02DF:q <= 8'h75;
            12'h02E0:q <= 8'h62;
            12'h02E1:q <= 8'h66;
            12'h02E2:q <= 8'hFF;
            12'h02E3:q <= 8'h18;
            12'h02E4:q <= 8'h6B;
            12'h02E5:q <= 8'h38;
            12'h02E6:q <= 8'hFF;
            12'h02E7:q <= 8'h00;
            12'h02E8:q <= 8'h0F;
            12'h02E9:q <= 8'h2D;
            12'h02EA:q <= 8'hFF;
            12'h02EB:q <= 8'h65;
            12'h02EC:q <= 8'h4F;
            12'h02ED:q <= 8'h0A;
            12'h02EE:q <= 8'hFF;
            12'h02EF:q <= 8'h13;
            12'h02F0:q <= 8'h03;
            12'h02F1:q <= 8'h01;
            12'h02F2:q <= 8'hFF;
            12'h02F3:q <= 8'h07;
            12'h02F4:q <= 8'h61;
            12'h02F5:q <= 8'h6C;
            12'h02F6:q <= 8'hFF;
            12'h02F7:q <= 8'h2C;
            12'h02F8:q <= 8'h21;
            12'h02F9:q <= 8'h4B;
            12'h02FA:q <= 8'hFF;
            12'h02FB:q <= 8'h58;
            12'h02FC:q <= 8'h55;
            12'h02FD:q <= 8'h6E;
            12'h02FE:q <= 8'hFF;
            12'h02FF:q <= 8'h3A;
            12'h0300:q <= 8'h36;
            12'h0301:q <= 8'h2F;
            12'h0302:q <= 8'hFF;
            12'h0303:q <= 8'h51;
            12'h0304:q <= 8'h40;
            12'h0305:q <= 8'h73;
            12'h0306:q <= 8'hFF;
            12'h0307:q <= 8'h24;
            12'h0308:q <= 8'h10;
            12'h0309:q <= 8'h6A;
            12'h030A:q <= 8'hFF;
            12'h030B:q <= 8'h22;
            12'h030C:q <= 8'h3E;
            12'h030D:q <= 8'h29;
            12'h030E:q <= 8'hFF;
            12'h030F:q <= 8'h01;
            12'h0310:q <= 8'h0C;
            12'h0311:q <= 8'h31;
            12'h0312:q <= 8'hFF;
            12'h0313:q <= 8'h1B;
            12'h0314:q <= 8'h66;
            12'h0315:q <= 8'h54;
            12'h0316:q <= 8'hFF;
            12'h0317:q <= 8'h4D;
            12'h0318:q <= 8'h68;
            12'h0319:q <= 8'h44;
            12'h031A:q <= 8'hFF;
            12'h031B:q <= 8'h1C;
            12'h031C:q <= 8'h51;
            12'h031D:q <= 8'h10;
            12'h031E:q <= 8'hFF;
            12'h031F:q <= 8'h30;
            12'h0320:q <= 8'h6C;
            12'h0321:q <= 8'h12;
            12'h0322:q <= 8'hFF;
            12'h0323:q <= 8'h21;
            12'h0324:q <= 8'h2A;
            12'h0325:q <= 8'h1F;
            12'h0326:q <= 8'hFF;
            12'h0327:q <= 8'h1A;
            12'h0328:q <= 8'h1D;
            12'h0329:q <= 8'h10;
            12'h032A:q <= 8'h06;
            12'h032B:q <= 8'h16;
            12'h032C:q <= 8'h0A;
            12'h032D:q <= 8'h02;
            12'h032E:q <= 8'h0F;
            12'h032F:q <= 8'h0D;
            12'h0330:q <= 8'h13;
            12'h0331:q <= 8'h03;
            12'h0332:q <= 8'h0C;
            12'h0333:q <= 8'hFF;
            12'h0334:q <= 8'h08;
            12'h0335:q <= 8'h0B;
            12'h0336:q <= 8'h13;
            12'h0337:q <= 8'h0C;
            12'h0338:q <= 8'h06;
            12'h0339:q <= 8'h11;
            12'h033A:q <= 8'h1C;
            12'h033B:q <= 8'h19;
            12'h033C:q <= 8'h01;
            12'h033D:q <= 8'h12;
            12'h033E:q <= 8'h06;
            12'h033F:q <= 8'h05;
            12'h0340:q <= 8'hFF;
            12'h0341:q <= 8'h17;
            12'h0342:q <= 8'h09;
            12'h0343:q <= 8'h04;
            12'h0344:q <= 8'h12;
            12'h0345:q <= 8'h07;
            12'h0346:q <= 8'h18;
            12'h0347:q <= 8'h00;
            12'h0348:q <= 8'h0E;
            12'h0349:q <= 8'h09;
            12'h034A:q <= 8'h1A;
            12'h034B:q <= 8'h0F;
            12'h034C:q <= 8'h0B;
            12'h034D:q <= 8'hFF;
            12'h034E:q <= 8'h07;
            12'h034F:q <= 8'h03;
            12'h0350:q <= 8'h19;
            12'h0351:q <= 8'h1B;
            12'h0352:q <= 8'h17;
            12'h0353:q <= 8'h15;
            12'h0354:q <= 8'h10;
            12'h0355:q <= 8'h05;
            12'h0356:q <= 8'h00;
            12'h0357:q <= 8'h0A;
            12'h0358:q <= 8'h16;
            12'h0359:q <= 8'h14;
            12'h035A:q <= 8'hFF;
            12'h035B:q <= 8'h14;
            12'h035C:q <= 8'h01;
            12'h035D:q <= 8'h0F;
            12'h035E:q <= 8'h18;
            12'h035F:q <= 8'h13;
            12'h0360:q <= 8'h1A;
            12'h0361:q <= 8'h0D;
            12'h0362:q <= 8'h01;
            12'h0363:q <= 8'h15;
            12'h0364:q <= 8'h1D;
            12'h0365:q <= 8'h02;
            12'h0366:q <= 8'h10;
            12'h0367:q <= 8'hFF;
            12'h0368:q <= 8'h05;
            12'h0369:q <= 8'h0C;
            12'h036A:q <= 8'h08;
            12'h036B:q <= 8'hFF;
            12'h036C:q <= 8'h02;
            12'h036D:q <= 8'h14;
            12'h036E:q <= 8'h17;
            12'h036F:q <= 8'hFF;
            12'h0370:q <= 8'h15;
            12'h0371:q <= 8'h0B;
            12'h0372:q <= 8'h19;
            12'h0373:q <= 8'hFF;
            12'h0374:q <= 8'h0A;
            12'h0375:q <= 8'h1D;
            12'h0376:q <= 8'h0E;
            12'h0377:q <= 8'hFF;
            12'h0378:q <= 8'h16;
            12'h0379:q <= 8'h03;
            12'h037A:q <= 8'h1C;
            12'h037B:q <= 8'hFF;
            12'h037C:q <= 8'h00;
            12'h037D:q <= 8'h12;
            12'h037E:q <= 8'h18;
            12'h037F:q <= 8'hFF;
            12'h0380:q <= 8'h0E;
            12'h0381:q <= 8'h09;
            12'h0382:q <= 8'h07;
            12'h0383:q <= 8'hFF;
            12'h0384:q <= 8'h0D;
            12'h0385:q <= 8'h1B;
            12'h0386:q <= 8'h04;
            12'h0387:q <= 8'hFF;
            12'h0388:q <= 8'h1C;
            12'h0389:q <= 8'h08;
            12'h038A:q <= 8'h1B;
            12'h038B:q <= 8'hFF;
            12'h038C:q <= 8'h11;
            12'h038D:q <= 8'h04;
            12'h038E:q <= 8'h11;
            12'h038F:q <= 8'hFF;
            12'h0390:q <= 8'h5D;
            12'h0391:q <= 8'h2A;
            12'h0392:q <= 8'h30;
            12'h0393:q <= 8'h53;
            12'h0394:q <= 8'h2E;
            12'h0395:q <= 8'h0C;
            12'h0396:q <= 8'h0D;
            12'h0397:q <= 8'h00;
            12'h0398:q <= 8'h17;
            12'h0399:q <= 8'h47;
            12'h039A:q <= 8'h22;
            12'h039B:q <= 8'h00;
            12'h039C:q <= 8'hFF;
            12'h039D:q <= 8'h68;
            12'h039E:q <= 8'h43;
            12'h039F:q <= 8'h46;
            12'h03A0:q <= 8'h03;
            12'h03A1:q <= 8'h54;
            12'h03A2:q <= 8'h6A;
            12'h03A3:q <= 8'h14;
            12'h03A4:q <= 8'h32;
            12'h03A5:q <= 8'h5E;
            12'h03A6:q <= 8'h49;
            12'h03A7:q <= 8'h1B;
            12'h03A8:q <= 8'h1D;
            12'h03A9:q <= 8'hFF;
            12'h03AA:q <= 8'h5F;
            12'h03AB:q <= 8'h6B;
            12'h03AC:q <= 8'h3A;
            12'h03AD:q <= 8'h16;
            12'h03AE:q <= 8'h50;
            12'h03AF:q <= 8'h25;
            12'h03B0:q <= 8'h09;
            12'h03B1:q <= 8'h3A;
            12'h03B2:q <= 8'h30;
            12'h03B3:q <= 8'h48;
            12'h03B4:q <= 8'h0C;
            12'h03B5:q <= 8'h2D;
            12'h03B6:q <= 8'hFF;
            12'h03B7:q <= 8'h5A;
            12'h03B8:q <= 8'h32;
            12'h03B9:q <= 8'h4F;
            12'h03BA:q <= 8'h61;
            12'h03BB:q <= 8'h31;
            12'h03BC:q <= 8'h69;
            12'h03BD:q <= 8'h1E;
            12'h03BE:q <= 8'h18;
            12'h03BF:q <= 8'h42;
            12'h03C0:q <= 8'h5B;
            12'h03C1:q <= 8'h4C;
            12'h03C2:q <= 8'h33;
            12'h03C3:q <= 8'hFF;
            12'h03C4:q <= 8'h1D;
            12'h03C5:q <= 8'h27;
            12'h03C6:q <= 8'h44;
            12'h03C7:q <= 8'h29;
            12'h03C8:q <= 8'h1A;
            12'h03C9:q <= 8'h3E;
            12'h03CA:q <= 8'h64;
            12'h03CB:q <= 8'h58;
            12'h03CC:q <= 8'h05;
            12'h03CD:q <= 8'h40;
            12'h03CE:q <= 8'h18;
            12'h03CF:q <= 8'h11;
            12'h03D0:q <= 8'hFF;
            12'h03D1:q <= 8'h41;
            12'h03D2:q <= 8'h05;
            12'h03D3:q <= 8'h14;
            12'h03D4:q <= 8'h18;
            12'h03D5:q <= 8'h29;
            12'h03D6:q <= 8'h53;
            12'h03D7:q <= 8'h04;
            12'h03D8:q <= 8'h40;
            12'h03D9:q <= 8'h6A;
            12'h03DA:q <= 8'h3C;
            12'h03DB:q <= 8'h66;
            12'h03DC:q <= 8'h5C;
            12'h03DD:q <= 8'hFF;
            12'h03DE:q <= 8'h55;
            12'h03DF:q <= 8'h23;
            12'h03E0:q <= 8'h13;
            12'h03E1:q <= 8'h3E;
            12'h03E2:q <= 8'h1C;
            12'h03E3:q <= 8'h5A;
            12'h03E4:q <= 8'h02;
            12'h03E5:q <= 8'h1F;
            12'h03E6:q <= 8'h36;
            12'h03E7:q <= 8'h1E;
            12'h03E8:q <= 8'h59;
            12'h03E9:q <= 8'h2F;
            12'h03EA:q <= 8'hFF;
            12'h03EB:q <= 8'h12;
            12'h03EC:q <= 8'h38;
            12'h03ED:q <= 8'h0D;
            12'h03EE:q <= 8'h50;
            12'h03EF:q <= 8'h68;
            12'h03F0:q <= 8'h2C;
            12'h03F1:q <= 8'h62;
            12'h03F2:q <= 8'h28;
            12'h03F3:q <= 8'h6B;
            12'h03F4:q <= 8'h45;
            12'h03F5:q <= 8'h15;
            12'h03F6:q <= 8'h50;
            12'h03F7:q <= 8'hFF;
            12'h03F8:q <= 8'h1A;
            12'h03F9:q <= 8'h49;
            12'h03FA:q <= 8'h1C;
            12'h03FB:q <= 8'h37;
            12'h03FC:q <= 8'h11;
            12'h03FD:q <= 8'h46;
            12'h03FE:q <= 8'h38;
            12'h03FF:q <= 8'h26;
            12'h0400:q <= 8'h13;
            12'h0401:q <= 8'h08;
            12'h0402:q <= 8'h43;
            12'h0403:q <= 8'h0D;
            12'h0404:q <= 8'hFF;
            12'h0405:q <= 8'h17;
            12'h0406:q <= 8'h6A;
            12'h0407:q <= 8'h36;
            12'h0408:q <= 8'h3B;
            12'h0409:q <= 8'h12;
            12'h040A:q <= 8'h21;
            12'h040B:q <= 8'h34;
            12'h040C:q <= 8'h5C;
            12'h040D:q <= 8'h58;
            12'h040E:q <= 8'h24;
            12'h040F:q <= 8'h07;
            12'h0410:q <= 8'h20;
            12'h0411:q <= 8'hFF;
            12'h0412:q <= 8'h4E;
            12'h0413:q <= 8'h09;
            12'h0414:q <= 8'h59;
            12'h0415:q <= 8'h06;
            12'h0416:q <= 8'h22;
            12'h0417:q <= 8'h17;
            12'h0418:q <= 8'h5F;
            12'h0419:q <= 8'h55;
            12'h041A:q <= 8'h53;
            12'h041B:q <= 8'h51;
            12'h041C:q <= 8'h56;
            12'h041D:q <= 8'h3A;
            12'h041E:q <= 8'hFF;
            12'h041F:q <= 8'h3D;
            12'h0420:q <= 8'h25;
            12'h0421:q <= 8'h31;
            12'h0422:q <= 8'h2D;
            12'h0423:q <= 8'h3C;
            12'h0424:q <= 8'h13;
            12'h0425:q <= 8'h0A;
            12'h0426:q <= 8'h47;
            12'h0427:q <= 8'h02;
            12'h0428:q <= 8'h2B;
            12'h0429:q <= 8'h1F;
            12'h042A:q <= 8'h27;
            12'h042B:q <= 8'hFF;
            12'h042C:q <= 8'h42;
            12'h042D:q <= 8'h0B;
            12'h042E:q <= 8'h39;
            12'h042F:q <= 8'h34;
            12'h0430:q <= 8'h4A;
            12'h0431:q <= 8'h16;
            12'h0432:q <= 8'h3B;
            12'h0433:q <= 8'h08;
            12'h0434:q <= 8'h4A;
            12'h0435:q <= 8'h26;
            12'h0436:q <= 8'h4F;
            12'h0437:q <= 8'h03;
            12'h0438:q <= 8'hFF;
            12'h0439:q <= 8'h5E;
            12'h043A:q <= 8'h33;
            12'h043B:q <= 8'h26;
            12'h043C:q <= 8'h67;
            12'h043D:q <= 8'h27;
            12'h043E:q <= 8'h4E;
            12'h043F:q <= 8'h36;
            12'h0440:q <= 8'h2D;
            12'h0441:q <= 8'h14;
            12'h0442:q <= 8'h04;
            12'h0443:q <= 8'h2A;
            12'h0444:q <= 8'h23;
            12'h0445:q <= 8'hFF;
            12'h0446:q <= 8'h2F;
            12'h0447:q <= 8'h0E;
            12'h0448:q <= 8'h56;
            12'h0449:q <= 8'h15;
            12'h044A:q <= 8'h5B;
            12'h044B:q <= 8'h05;
            12'h044C:q <= 8'h63;
            12'h044D:q <= 8'h66;
            12'h044E:q <= 8'h5F;
            12'h044F:q <= 8'h4E;
            12'h0450:q <= 8'h0F;
            12'h0451:q <= 8'h3D;
            12'h0452:q <= 8'hFF;
            12'h0453:q <= 8'h4C;
            12'h0454:q <= 8'h22;
            12'h0455:q <= 8'h20;
            12'h0456:q <= 8'h10;
            12'h0457:q <= 8'h6B;
            12'h0458:q <= 8'h24;
            12'h0459:q <= 8'h65;
            12'h045A:q <= 8'h56;
            12'h045B:q <= 8'h0B;
            12'h045C:q <= 8'h5A;
            12'h045D:q <= 8'h64;
            12'h045E:q <= 8'h2C;
            12'h045F:q <= 8'hFF;
            12'h0460:q <= 8'h63;
            12'h0461:q <= 8'h1B;
            12'h0462:q <= 8'h2C;
            12'h0463:q <= 8'h04;
            12'h0464:q <= 8'h39;
            12'h0465:q <= 8'h19;
            12'h0466:q <= 8'h42;
            12'h0467:q <= 8'h41;
            12'h0468:q <= 8'h28;
            12'h0469:q <= 8'h5D;
            12'h046A:q <= 8'h16;
            12'h046B:q <= 8'h44;
            12'h046C:q <= 8'hFF;
            12'h046D:q <= 8'h21;
            12'h046E:q <= 8'h57;
            12'h046F:q <= 8'h01;
            12'h0470:q <= 8'h24;
            12'h0471:q <= 8'h0B;
            12'h0472:q <= 8'h10;
            12'h0473:q <= 8'h35;
            12'h0474:q <= 8'h06;
            12'h0475:q <= 8'h63;
            12'h0476:q <= 8'h06;
            12'h0477:q <= 8'h62;
            12'h0478:q <= 8'h65;
            12'h0479:q <= 8'hFF;
            12'h047A:q <= 8'h0A;
            12'h047B:q <= 8'h2B;
            12'h047C:q <= 8'h4B;
            12'h047D:q <= 8'h1E;
            12'h047E:q <= 8'h4F;
            12'h047F:q <= 8'h48;
            12'h0480:q <= 8'h2A;
            12'h0481:q <= 8'h20;
            12'h0482:q <= 8'h37;
            12'h0483:q <= 8'h35;
            12'h0484:q <= 8'h55;
            12'h0485:q <= 8'h3F;
            12'h0486:q <= 8'hFF;
            12'h0487:q <= 8'h45;
            12'h0488:q <= 8'h19;
            12'h0489:q <= 8'h51;
            12'h048A:q <= 8'h40;
            12'h048B:q <= 8'h3F;
            12'h048C:q <= 8'h37;
            12'h048D:q <= 8'h2F;
            12'h048E:q <= 8'h01;
            12'h048F:q <= 8'h29;
            12'h0490:q <= 8'h09;
            12'h0491:q <= 8'h1A;
            12'h0492:q <= 8'h46;
            12'h0493:q <= 8'hFF;
            12'h0494:q <= 8'h08;
            12'h0495:q <= 8'h66;
            12'h0496:q <= 8'h52;
            12'h0497:q <= 8'h54;
            12'h0498:q <= 8'h5E;
            12'h0499:q <= 8'h49;
            12'h049A:q <= 8'h52;
            12'h049B:q <= 8'h3D;
            12'h049C:q <= 8'h54;
            12'h049D:q <= 8'h31;
            12'h049E:q <= 8'h61;
            12'h049F:q <= 8'h57;
            12'h04A0:q <= 8'hFF;
            12'h04A1:q <= 8'h65;
            12'h04A2:q <= 8'h4D;
            12'h04A3:q <= 8'h48;
            12'h04A4:q <= 8'h0C;
            12'h04A5:q <= 8'h67;
            12'h04A6:q <= 8'h61;
            12'h04A7:q <= 8'h30;
            12'h04A8:q <= 8'h23;
            12'h04A9:q <= 8'h67;
            12'h04AA:q <= 8'h10;
            12'h04AB:q <= 8'h0A;
            12'h04AC:q <= 8'h12;
            12'h04AD:q <= 8'hFF;
            12'h04AE:q <= 8'h3F;
            12'h04AF:q <= 8'h0F;
            12'h04B0:q <= 8'h28;
            12'h04B1:q <= 8'h35;
            12'h04B2:q <= 8'h15;
            12'h04B3:q <= 8'h5D;
            12'h04B4:q <= 8'h1B;
            12'h04B5:q <= 8'h51;
            12'h04B6:q <= 8'h69;
            12'h04B7:q <= 8'h68;
            12'h04B8:q <= 8'h39;
            12'h04B9:q <= 8'h4D;
            12'h04BA:q <= 8'hFF;
            12'h04BB:q <= 8'h47;
            12'h04BC:q <= 8'h2E;
            12'h04BD:q <= 8'h11;
            12'h04BE:q <= 8'h60;
            12'h04BF:q <= 8'h03;
            12'h04C0:q <= 8'h59;
            12'h04C1:q <= 8'h0F;
            12'h04C2:q <= 8'h1D;
            12'h04C3:q <= 8'h32;
            12'h04C4:q <= 8'h52;
            12'h04C5:q <= 8'h3E;
            12'h04C6:q <= 8'h01;
            12'h04C7:q <= 8'hFF;
            12'h04C8:q <= 8'h07;
            12'h04C9:q <= 8'h4C;
            12'h04CA:q <= 8'h19;
            12'h04CB:q <= 8'hFF;
            12'h04CC:q <= 8'h5C;
            12'h04CD:q <= 8'h2B;
            12'h04CE:q <= 8'h38;
            12'h04CF:q <= 8'hFF;
            12'h04D0:q <= 8'h58;
            12'h04D1:q <= 8'h60;
            12'h04D2:q <= 8'h0E;
            12'h04D3:q <= 8'hFF;
            12'h04D4:q <= 8'h1F;
            12'h04D5:q <= 8'h0E;
            12'h04D6:q <= 8'h34;
            12'h04D7:q <= 8'hFF;
            12'h04D8:q <= 8'h02;
            12'h04D9:q <= 8'h57;
            12'h04DA:q <= 8'h60;
            12'h04DB:q <= 8'hFF;
            12'h04DC:q <= 8'h64;
            12'h04DD:q <= 8'h4B;
            12'h04DE:q <= 8'h41;
            12'h04DF:q <= 8'hFF;
            12'h04E0:q <= 8'h5B;
            12'h04E1:q <= 8'h43;
            12'h04E2:q <= 8'h4B;
            12'h04E3:q <= 8'hFF;
            12'h04E4:q <= 8'h4A;
            12'h04E5:q <= 8'h4D;
            12'h04E6:q <= 8'h21;
            12'h04E7:q <= 8'hFF;
            12'h04E8:q <= 8'h00;
            12'h04E9:q <= 8'h07;
            12'h04EA:q <= 8'h2E;
            12'h04EB:q <= 8'hFF;
            12'h04EC:q <= 8'h3C;
            12'h04ED:q <= 8'h44;
            12'h04EE:q <= 8'h25;
            12'h04EF:q <= 8'hFF;
            12'h04F0:q <= 8'h69;
            12'h04F1:q <= 8'h33;
            12'h04F2:q <= 8'h1C;
            12'h04F3:q <= 8'hFF;
            12'h04F4:q <= 8'h62;
            12'h04F5:q <= 8'h45;
            12'h04F6:q <= 8'h3B;
            12'h04F7:q <= 8'hFF;
            12'h04F8:q <= 8'h5B;
            12'h04F9:q <= 8'h43;
            12'h04FA:q <= 8'h58;
            12'h04FB:q <= 8'hFF;
            12'h04FC:q <= 8'h31;
            12'h04FD:q <= 8'h2D;
            12'h04FE:q <= 8'h27;
            12'h04FF:q <= 8'hFF;
            12'h0500:q <= 8'h20;
            12'h0501:q <= 8'h4C;
            12'h0502:q <= 8'h36;
            12'h0503:q <= 8'hFF;
            12'h0504:q <= 8'h64;
            12'h0505:q <= 8'h1B;
            12'h0506:q <= 8'h52;
            12'h0507:q <= 8'hFF;
            12'h0508:q <= 8'h63;
            12'h0509:q <= 8'h3E;
            12'h050A:q <= 8'h02;
            12'h050B:q <= 8'hFF;
            12'h050C:q <= 8'h30;
            12'h050D:q <= 8'h6B;
            12'h050E:q <= 8'h3C;
            12'h050F:q <= 8'hFF;
            12'h0510:q <= 8'h44;
            12'h0511:q <= 8'h46;
            12'h0512:q <= 8'h0B;
            12'h0513:q <= 8'hFF;
            12'h0514:q <= 8'h60;
            12'h0515:q <= 8'h09;
            12'h0516:q <= 8'h49;
            12'h0517:q <= 8'hFF;
            12'h0518:q <= 8'h66;
            12'h0519:q <= 8'h33;
            12'h051A:q <= 8'h06;
            12'h051B:q <= 8'hFF;
            12'h051C:q <= 8'h01;
            12'h051D:q <= 8'h5E;
            12'h051E:q <= 8'h40;
            12'h051F:q <= 8'hFF;
            12'h0520:q <= 8'h08;
            12'h0521:q <= 8'h0C;
            12'h0522:q <= 8'h3D;
            12'h0523:q <= 8'hFF;
            12'h0524:q <= 8'h65;
            12'h0525:q <= 8'h3A;
            12'h0526:q <= 8'h0E;
            12'h0527:q <= 8'hFF;
            12'h0528:q <= 8'h15;
            12'h0529:q <= 8'h24;
            12'h052A:q <= 8'h4B;
            12'h052B:q <= 8'hFF;
            12'h052C:q <= 8'h45;
            12'h052D:q <= 8'h18;
            12'h052E:q <= 8'h03;
            12'h052F:q <= 8'hFF;
            12'h0530:q <= 8'h29;
            12'h0531:q <= 8'h28;
            12'h0532:q <= 8'h1C;
            12'h0533:q <= 8'hFF;
            12'h0534:q <= 8'h41;
            12'h0535:q <= 8'h3B;
            12'h0536:q <= 8'h1E;
            12'h0537:q <= 8'hFF;
            12'h0538:q <= 8'h54;
            12'h0539:q <= 8'h32;
            12'h053A:q <= 8'h38;
            12'h053B:q <= 8'hFF;
            12'h053C:q <= 8'h1A;
            12'h053D:q <= 8'h4A;
            12'h053E:q <= 8'h1F;
            12'h053F:q <= 8'hFF;
            12'h0540:q <= 8'h67;
            12'h0541:q <= 8'h47;
            12'h0542:q <= 8'h5C;
            12'h0543:q <= 8'hFF;
            12'h0544:q <= 8'h48;
            12'h0545:q <= 8'h5A;
            12'h0546:q <= 8'h59;
            12'h0547:q <= 8'hFF;
            12'h0548:q <= 8'h19;
            12'h0549:q <= 8'h61;
            12'h054A:q <= 8'h16;
            12'h054B:q <= 8'hFF;
            12'h054C:q <= 8'h37;
            12'h054D:q <= 8'h0F;
            12'h054E:q <= 8'h22;
            12'h054F:q <= 8'hFF;
            12'h0550:q <= 8'h2E;
            12'h0551:q <= 8'h2A;
            12'h0552:q <= 8'h42;
            12'h0553:q <= 8'hFF;
            12'h0554:q <= 8'h10;
            12'h0555:q <= 8'h14;
            12'h0556:q <= 8'h11;
            12'h0557:q <= 8'hFF;
            12'h0558:q <= 8'h5F;
            12'h0559:q <= 8'h56;
            12'h055A:q <= 8'h0D;
            12'h055B:q <= 8'hFF;
            12'h055C:q <= 8'h50;
            12'h055D:q <= 8'h62;
            12'h055E:q <= 8'h07;
            12'h055F:q <= 8'hFF;
            12'h0560:q <= 8'h68;
            12'h0561:q <= 8'h35;
            12'h0562:q <= 8'h26;
            12'h0563:q <= 8'hFF;
            12'h0564:q <= 8'h6A;
            12'h0565:q <= 8'h51;
            12'h0566:q <= 8'h12;
            12'h0567:q <= 8'hFF;
            12'h0568:q <= 8'h69;
            12'h0569:q <= 8'h39;
            12'h056A:q <= 8'h1D;
            12'h056B:q <= 8'hFF;
            12'h056C:q <= 8'h55;
            12'h056D:q <= 8'h25;
            12'h056E:q <= 8'h17;
            12'h056F:q <= 8'hFF;
            12'h0570:q <= 8'h05;
            12'h0571:q <= 8'h57;
            12'h0572:q <= 8'h3F;
            12'h0573:q <= 8'hFF;
            12'h0574:q <= 8'h53;
            12'h0575:q <= 8'h23;
            12'h0576:q <= 8'h0A;
            12'h0577:q <= 8'hFF;
            12'h0578:q <= 8'h13;
            12'h0579:q <= 8'h2F;
            12'h057A:q <= 8'h2B;
            12'h057B:q <= 8'hFF;
            12'h057C:q <= 8'h2C;
            12'h057D:q <= 8'h21;
            12'h057E:q <= 8'h34;
            12'h057F:q <= 8'hFF;
            12'h0580:q <= 8'h4D;
            12'h0581:q <= 8'h5D;
            12'h0582:q <= 8'h4E;
            12'h0583:q <= 8'hFF;
            12'h0584:q <= 8'h00;
            12'h0585:q <= 8'h4F;
            12'h0586:q <= 8'h04;
            12'h0587:q <= 8'hFF;
            12'h0588:q <= 8'h07;
            12'h0589:q <= 8'h0C;
            12'h058A:q <= 8'h02;
            12'h058B:q <= 8'h10;
            12'h058C:q <= 8'h18;
            12'h058D:q <= 8'h19;
            12'h058E:q <= 8'h0E;
            12'h058F:q <= 8'h0C;
            12'h0590:q <= 8'h15;
            12'h0591:q <= 8'h0A;
            12'h0592:q <= 8'h09;
            12'h0593:q <= 8'h10;
            12'h0594:q <= 8'hFF;
            12'h0595:q <= 8'h1A;
            12'h0596:q <= 8'h0B;
            12'h0597:q <= 8'h15;
            12'h0598:q <= 8'h0A;
            12'h0599:q <= 8'h1A;
            12'h059A:q <= 8'h01;
            12'h059B:q <= 8'h13;
            12'h059C:q <= 8'h0D;
            12'h059D:q <= 8'h14;
            12'h059E:q <= 8'h03;
            12'h059F:q <= 8'h0F;
            12'h05A0:q <= 8'h18;
            12'h05A1:q <= 8'hFF;
            12'h05A2:q <= 8'h17;
            12'h05A3:q <= 8'h0F;
            12'h05A4:q <= 8'h03;
            12'h05A5:q <= 8'h16;
            12'h05A6:q <= 8'h06;
            12'h05A7:q <= 8'h10;
            12'h05A8:q <= 8'h14;
            12'h05A9:q <= 8'h03;
            12'h05AA:q <= 8'h08;
            12'h05AB:q <= 8'h0C;
            12'h05AC:q <= 8'h16;
            12'h05AD:q <= 8'h0E;
            12'h05AE:q <= 8'hFF;
            12'h05AF:q <= 8'h04;
            12'h05B0:q <= 8'h01;
            12'h05B1:q <= 8'h11;
            12'h05B2:q <= 8'h06;
            12'h05B3:q <= 8'h07;
            12'h05B4:q <= 8'h12;
            12'h05B5:q <= 8'h17;
            12'h05B6:q <= 8'h08;
            12'h05B7:q <= 8'h00;
            12'h05B8:q <= 8'h19;
            12'h05B9:q <= 8'h11;
            12'h05BA:q <= 8'h0D;
            12'h05BB:q <= 8'hFF;
            12'h05BC:q <= 8'h08;
            12'h05BD:q <= 8'h18;
            12'h05BE:q <= 8'h14;
            12'h05BF:q <= 8'h13;
            12'h05C0:q <= 8'h15;
            12'h05C1:q <= 8'h00;
            12'h05C2:q <= 8'h05;
            12'h05C3:q <= 8'h16;
            12'h05C4:q <= 8'h0B;
            12'h05C5:q <= 8'h05;
            12'h05C6:q <= 8'h06;
            12'h05C7:q <= 8'h1A;
            12'h05C8:q <= 8'hFF;
            12'h05C9:q <= 8'h00;
            12'h05CA:q <= 8'h0E;
            12'h05CB:q <= 8'h09;
            12'h05CC:q <= 8'h0D;
            12'h05CD:q <= 8'h02;
            12'h05CE:q <= 8'h0F;
            12'h05CF:q <= 8'h0B;
            12'h05D0:q <= 8'h0A;
            12'h05D1:q <= 8'h07;
            12'h05D2:q <= 8'h12;
            12'h05D3:q <= 8'h17;
            12'h05D4:q <= 8'h02;
            12'h05D5:q <= 8'hFF;
            12'h05D6:q <= 8'h05;
            12'h05D7:q <= 8'h11;
            12'h05D8:q <= 8'h04;
            12'h05D9:q <= 8'hFF;
            12'h05DA:q <= 8'h12;
            12'h05DB:q <= 8'h09;
            12'h05DC:q <= 8'h13;
            12'h05DD:q <= 8'hFF;
            12'h05DE:q <= 8'h19;
            12'h05DF:q <= 8'h04;
            12'h05E0:q <= 8'h01;
            12'h05E1:q <= 8'hFF;
            12'h05E2:q <= 8'h1A;
            12'h05E3:q <= 8'h0C;
            12'h05E4:q <= 8'h08;
            12'h05E5:q <= 8'hFF;
            12'h05E6:q <= 8'h09;
            12'h05E7:q <= 8'h15;
            12'h05E8:q <= 8'h11;
            12'h05E9:q <= 8'hFF;
            12'h05EA:q <= 8'h0F;
            12'h05EB:q <= 8'h12;
            12'h05EC:q <= 8'h0D;
            12'h05ED:q <= 8'hFF;
            12'h05EE:q <= 8'h10;
            12'h05EF:q <= 8'h07;
            12'h05F0:q <= 8'h05;
            12'h05F1:q <= 8'hFF;
            12'h05F2:q <= 8'h02;
            12'h05F3:q <= 8'h16;
            12'h05F4:q <= 8'h06;
            12'h05F5:q <= 8'hFF;
            12'h05F6:q <= 8'h01;
            12'h05F7:q <= 8'h18;
            12'h05F8:q <= 8'h03;
            12'h05F9:q <= 8'hFF;
            12'h05FA:q <= 8'h14;
            12'h05FB:q <= 8'h0B;
            12'h05FC:q <= 8'h17;
            12'h05FD:q <= 8'hFF;
            12'h05FE:q <= 8'h04;
            12'h05FF:q <= 8'h19;
            12'h0600:q <= 8'h13;
            12'h0601:q <= 8'hFF;
            12'h0602:q <= 8'h0A;
            12'h0603:q <= 8'h00;
            12'h0604:q <= 8'h0E;
            12'h0605:q <= 8'hFF;
            12'h0606:q <= 8'h36;
            12'h0607:q <= 8'h30;
            12'h0608:q <= 8'h52;
            12'h0609:q <= 8'h15;
            12'h060A:q <= 8'h59;
            12'h060B:q <= 8'h31;
            12'h060C:q <= 8'h0E;
            12'h060D:q <= 8'h2F;
            12'h060E:q <= 8'hFF;
            12'h060F:q <= 8'h37;
            12'h0610:q <= 8'h3F;
            12'h0611:q <= 8'h2D;
            12'h0612:q <= 8'h0A;
            12'h0613:q <= 8'h32;
            12'h0614:q <= 8'h3F;
            12'h0615:q <= 8'h46;
            12'h0616:q <= 8'h33;
            12'h0617:q <= 8'hFF;
            12'h0618:q <= 8'h38;
            12'h0619:q <= 8'h47;
            12'h061A:q <= 8'h03;
            12'h061B:q <= 8'h1A;
            12'h061C:q <= 8'h13;
            12'h061D:q <= 8'h50;
            12'h061E:q <= 8'h48;
            12'h061F:q <= 8'h4F;
            12'h0620:q <= 8'hFF;
            12'h0621:q <= 8'h39;
            12'h0622:q <= 8'h33;
            12'h0623:q <= 8'h36;
            12'h0624:q <= 8'h17;
            12'h0625:q <= 8'h1F;
            12'h0626:q <= 8'h39;
            12'h0627:q <= 8'h05;
            12'h0628:q <= 8'h40;
            12'h0629:q <= 8'hFF;
            12'h062A:q <= 8'h3A;
            12'h062B:q <= 8'h0A;
            12'h062C:q <= 8'h07;
            12'h062D:q <= 8'h3A;
            12'h062E:q <= 8'h02;
            12'h062F:q <= 8'h18;
            12'h0630:q <= 8'h1F;
            12'h0631:q <= 8'h25;
            12'h0632:q <= 8'hFF;
            12'h0633:q <= 8'h3B;
            12'h0634:q <= 8'h31;
            12'h0635:q <= 8'h58;
            12'h0636:q <= 8'h1D;
            12'h0637:q <= 8'h2D;
            12'h0638:q <= 8'h34;
            12'h0639:q <= 8'h0A;
            12'h063A:q <= 8'h24;
            12'h063B:q <= 8'hFF;
            12'h063C:q <= 8'h3C;
            12'h063D:q <= 8'h38;
            12'h063E:q <= 8'h1D;
            12'h063F:q <= 8'h44;
            12'h0640:q <= 8'h03;
            12'h0641:q <= 8'h10;
            12'h0642:q <= 8'h36;
            12'h0643:q <= 8'h20;
            12'h0644:q <= 8'hFF;
            12'h0645:q <= 8'h3D;
            12'h0646:q <= 8'h42;
            12'h0647:q <= 8'h53;
            12'h0648:q <= 8'h4D;
            12'h0649:q <= 8'h2E;
            12'h064A:q <= 8'h58;
            12'h064B:q <= 8'h1B;
            12'h064C:q <= 8'h26;
            12'h064D:q <= 8'hFF;
            12'h064E:q <= 8'h3E;
            12'h064F:q <= 8'h15;
            12'h0650:q <= 8'h0B;
            12'h0651:q <= 8'h56;
            12'h0652:q <= 8'h36;
            12'h0653:q <= 8'h0D;
            12'h0654:q <= 8'h11;
            12'h0655:q <= 8'h2C;
            12'h0656:q <= 8'hFF;
            12'h0657:q <= 8'h3F;
            12'h0658:q <= 8'h43;
            12'h0659:q <= 8'h17;
            12'h065A:q <= 8'h4A;
            12'h065B:q <= 8'h04;
            12'h065C:q <= 8'h55;
            12'h065D:q <= 8'h4A;
            12'h065E:q <= 8'h52;
            12'h065F:q <= 8'hFF;
            12'h0660:q <= 8'h40;
            12'h0661:q <= 8'h25;
            12'h0662:q <= 8'h01;
            12'h0663:q <= 8'h35;
            12'h0664:q <= 8'h55;
            12'h0665:q <= 8'h26;
            12'h0666:q <= 8'h30;
            12'h0667:q <= 8'h01;
            12'h0668:q <= 8'hFF;
            12'h0669:q <= 8'h41;
            12'h066A:q <= 8'h14;
            12'h066B:q <= 8'h54;
            12'h066C:q <= 8'h57;
            12'h066D:q <= 8'h22;
            12'h066E:q <= 8'h32;
            12'h066F:q <= 8'h15;
            12'h0670:q <= 8'h10;
            12'h0671:q <= 8'hFF;
            12'h0672:q <= 8'h42;
            12'h0673:q <= 8'h32;
            12'h0674:q <= 8'h3E;
            12'h0675:q <= 8'h3C;
            12'h0676:q <= 8'h39;
            12'h0677:q <= 8'h3D;
            12'h0678:q <= 8'h22;
            12'h0679:q <= 8'h3E;
            12'h067A:q <= 8'hFF;
            12'h067B:q <= 8'h43;
            12'h067C:q <= 8'h46;
            12'h067D:q <= 8'h05;
            12'h067E:q <= 8'h50;
            12'h067F:q <= 8'h1B;
            12'h0680:q <= 8'h4E;
            12'h0681:q <= 8'h0F;
            12'h0682:q <= 8'h41;
            12'h0683:q <= 8'hFF;
            12'h0684:q <= 8'h44;
            12'h0685:q <= 8'h1D;
            12'h0686:q <= 8'h30;
            12'h0687:q <= 8'h4C;
            12'h0688:q <= 8'h12;
            12'h0689:q <= 8'h06;
            12'h068A:q <= 8'h2B;
            12'h068B:q <= 8'h23;
            12'h068C:q <= 8'hFF;
            12'h068D:q <= 8'h45;
            12'h068E:q <= 8'h0C;
            12'h068F:q <= 8'h13;
            12'h0690:q <= 8'h58;
            12'h0691:q <= 8'h42;
            12'h0692:q <= 8'h28;
            12'h0693:q <= 8'h21;
            12'h0694:q <= 8'h4E;
            12'h0695:q <= 8'hFF;
            12'h0696:q <= 8'h46;
            12'h0697:q <= 8'h02;
            12'h0698:q <= 8'h2A;
            12'h0699:q <= 8'h08;
            12'h069A:q <= 8'h0D;
            12'h069B:q <= 8'h03;
            12'h069C:q <= 8'h51;
            12'h069D:q <= 8'h21;
            12'h069E:q <= 8'hFF;
            12'h069F:q <= 8'h47;
            12'h06A0:q <= 8'h18;
            12'h06A1:q <= 8'h20;
            12'h06A2:q <= 8'h29;
            12'h06A3:q <= 8'h47;
            12'h06A4:q <= 8'h3B;
            12'h06A5:q <= 8'h41;
            12'h06A6:q <= 8'h34;
            12'h06A7:q <= 8'hFF;
            12'h06A8:q <= 8'h48;
            12'h06A9:q <= 8'h08;
            12'h06AA:q <= 8'h40;
            12'h06AB:q <= 8'h49;
            12'h06AC:q <= 8'h0E;
            12'h06AD:q <= 8'h1C;
            12'h06AE:q <= 8'h54;
            12'h06AF:q <= 8'h2D;
            12'h06B0:q <= 8'hFF;
            12'h06B1:q <= 8'h49;
            12'h06B2:q <= 8'h59;
            12'h06B3:q <= 8'h19;
            12'h06B4:q <= 8'h0B;
            12'h06B5:q <= 8'h14;
            12'h06B6:q <= 8'h2C;
            12'h06B7:q <= 8'h16;
            12'h06B8:q <= 8'h17;
            12'h06B9:q <= 8'hFF;
            12'h06BA:q <= 8'h4A;
            12'h06BB:q <= 8'h0B;
            12'h06BC:q <= 8'h46;
            12'h06BD:q <= 8'h28;
            12'h06BE:q <= 8'h2A;
            12'h06BF:q <= 8'h27;
            12'h06C0:q <= 8'h1E;
            12'h06C1:q <= 8'h01;
            12'h06C2:q <= 8'hFF;
            12'h06C3:q <= 8'h4B;
            12'h06C4:q <= 8'h06;
            12'h06C5:q <= 8'h2E;
            12'h06C6:q <= 8'h2B;
            12'h06C7:q <= 8'h09;
            12'h06C8:q <= 8'h24;
            12'h06C9:q <= 8'h33;
            12'h06CA:q <= 8'h3C;
            12'h06CB:q <= 8'hFF;
            12'h06CC:q <= 8'h4C;
            12'h06CD:q <= 8'h2D;
            12'h06CE:q <= 8'h4A;
            12'h06CF:q <= 8'h1E;
            12'h06D0:q <= 8'h45;
            12'h06D1:q <= 8'h23;
            12'h06D2:q <= 8'h4F;
            12'h06D3:q <= 8'h4B;
            12'h06D4:q <= 8'hFF;
            12'h06D5:q <= 8'h4D;
            12'h06D6:q <= 8'h3A;
            12'h06D7:q <= 8'h12;
            12'h06D8:q <= 8'h4B;
            12'h06D9:q <= 8'h0F;
            12'h06DA:q <= 8'h35;
            12'h06DB:q <= 8'h56;
            12'h06DC:q <= 8'h40;
            12'h06DD:q <= 8'hFF;
            12'h06DE:q <= 8'h4E;
            12'h06DF:q <= 8'h04;
            12'h06E0:q <= 8'h4D;
            12'h06E1:q <= 8'h05;
            12'h06E2:q <= 8'h19;
            12'h06E3:q <= 8'h42;
            12'h06E4:q <= 8'h47;
            12'h06E5:q <= 8'h09;
            12'h06E6:q <= 8'hFF;
            12'h06E7:q <= 8'h4F;
            12'h06E8:q <= 8'h2C;
            12'h06E9:q <= 8'h24;
            12'h06EA:q <= 8'h37;
            12'h06EB:q <= 8'h1C;
            12'h06EC:q <= 8'h20;
            12'h06ED:q <= 8'h12;
            12'h06EE:q <= 8'h57;
            12'h06EF:q <= 8'hFF;
            12'h06F0:q <= 8'h50;
            12'h06F1:q <= 8'h4C;
            12'h06F2:q <= 8'h39;
            12'h06F3:q <= 8'h27;
            12'h06F4:q <= 8'h00;
            12'h06F5:q <= 8'h2F;
            12'h06F6:q <= 8'h45;
            12'h06F7:q <= 8'h0C;
            12'h06F8:q <= 8'hFF;
            12'h06F9:q <= 8'h51;
            12'h06FA:q <= 8'h49;
            12'h06FB:q <= 8'h00;
            12'h06FC:q <= 8'h53;
            12'h06FD:q <= 8'h11;
            12'h06FE:q <= 8'h02;
            12'h06FF:q <= 8'h19;
            12'h0700:q <= 8'h2A;
            12'h0701:q <= 8'hFF;
            12'h0702:q <= 8'h52;
            12'h0703:q <= 8'h23;
            12'h0704:q <= 8'h47;
            12'h0705:q <= 8'h54;
            12'h0706:q <= 8'h07;
            12'h0707:q <= 8'h13;
            12'h0708:q <= 8'h4D;
            12'h0709:q <= 8'h38;
            12'h070A:q <= 8'hFF;
            12'h070B:q <= 8'h53;
            12'h070C:q <= 8'h55;
            12'h070D:q <= 8'h31;
            12'h070E:q <= 8'h3B;
            12'h070F:q <= 8'h3F;
            12'h0710:q <= 8'h4C;
            12'h0711:q <= 8'h1A;
            12'h0712:q <= 8'h3A;
            12'h0713:q <= 8'hFF;
            12'h0714:q <= 8'h54;
            12'h0715:q <= 8'h05;
            12'h0716:q <= 8'h0F;
            12'h0717:q <= 8'h38;
            12'h0718:q <= 8'h43;
            12'h0719:q <= 8'h08;
            12'h071A:q <= 8'h00;
            12'h071B:q <= 8'h37;
            12'h071C:q <= 8'hFF;
            12'h071D:q <= 8'h55;
            12'h071E:q <= 8'h56;
            12'h071F:q <= 8'h44;
            12'h0720:q <= 8'h16;
            12'h0721:q <= 8'h3D;
            12'h0722:q <= 8'h14;
            12'h0723:q <= 8'h25;
            12'h0724:q <= 8'h29;
            12'h0725:q <= 8'hFF;
            12'h0726:q <= 8'h56;
            12'h0727:q <= 8'h1C;
            12'h0728:q <= 8'h56;
            12'h0729:q <= 8'h06;
            12'h072A:q <= 8'h46;
            12'h072B:q <= 8'h0B;
            12'h072C:q <= 8'h59;
            12'h072D:q <= 8'h44;
            12'h072E:q <= 8'hFF;
            12'h072F:q <= 8'h57;
            12'h0730:q <= 8'h40;
            12'h0731:q <= 8'h55;
            12'h0732:q <= 8'h31;
            12'h0733:q <= 8'h0C;
            12'h0734:q <= 8'h2E;
            12'h0735:q <= 8'h04;
            12'h0736:q <= 8'h53;
            12'h0737:q <= 8'hFF;
            12'h0738:q <= 8'h58;
            12'h0739:q <= 8'h1B;
            12'h073A:q <= 8'h3F;
            12'h073B:q <= 8'h51;
            12'h073C:q <= 8'h48;
            12'h073D:q <= 8'h07;
            12'h073E:q <= 8'h52;
            12'h073F:q <= 8'h43;
            12'h0740:q <= 8'hFF;
            12'h0741:q <= 8'h59;
            12'h0742:q <= 8'h21;
            12'h0743:q <= 8'h3A;
            12'h0744:q <= 8'h30;
            12'h0745:q <= 8'h18;
            12'h0746:q <= 8'h3E;
            12'h0747:q <= 8'h1D;
            12'h0748:q <= 8'h49;
            12'h0749:q <= 8'hFF;
            12'h074A:q <= 8'h00;
            12'h074B:q <= 8'h4D;
            12'h074C:q <= 8'h23;
            12'h074D:q <= 8'hFF;
            12'h074E:q <= 8'h01;
            12'h074F:q <= 8'h26;
            12'h0750:q <= 8'h0A;
            12'h0751:q <= 8'hFF;
            12'h0752:q <= 8'h02;
            12'h0753:q <= 8'h13;
            12'h0754:q <= 8'h3C;
            12'h0755:q <= 8'hFF;
            12'h0756:q <= 8'h03;
            12'h0757:q <= 8'h48;
            12'h0758:q <= 8'h2C;
            12'h0759:q <= 8'hFF;
            12'h075A:q <= 8'h04;
            12'h075B:q <= 8'h35;
            12'h075C:q <= 8'h21;
            12'h075D:q <= 8'hFF;
            12'h075E:q <= 8'h05;
            12'h075F:q <= 8'h01;
            12'h0760:q <= 8'h4E;
            12'h0761:q <= 8'hFF;
            12'h0762:q <= 8'h06;
            12'h0763:q <= 8'h57;
            12'h0764:q <= 8'h38;
            12'h0765:q <= 8'hFF;
            12'h0766:q <= 8'h07;
            12'h0767:q <= 8'h44;
            12'h0768:q <= 8'h59;
            12'h0769:q <= 8'hFF;
            12'h076A:q <= 8'h08;
            12'h076B:q <= 8'h4E;
            12'h076C:q <= 8'h3B;
            12'h076D:q <= 8'hFF;
            12'h076E:q <= 8'h09;
            12'h076F:q <= 8'h17;
            12'h0770:q <= 8'h1C;
            12'h0771:q <= 8'hFF;
            12'h0772:q <= 8'h0A;
            12'h0773:q <= 8'h1F;
            12'h0774:q <= 8'h0D;
            12'h0775:q <= 8'hFF;
            12'h0776:q <= 8'h0B;
            12'h0777:q <= 8'h1E;
            12'h0778:q <= 8'h41;
            12'h0779:q <= 8'hFF;
            12'h077A:q <= 8'h0C;
            12'h077B:q <= 8'h27;
            12'h077C:q <= 8'h4F;
            12'h077D:q <= 8'hFF;
            12'h077E:q <= 8'h0D;
            12'h077F:q <= 8'h11;
            12'h0780:q <= 8'h43;
            12'h0781:q <= 8'hFF;
            12'h0782:q <= 8'h0E;
            12'h0783:q <= 8'h2F;
            12'h0784:q <= 8'h26;
            12'h0785:q <= 8'hFF;
            12'h0786:q <= 8'h0F;
            12'h0787:q <= 8'h24;
            12'h0788:q <= 8'h02;
            12'h0789:q <= 8'hFF;
            12'h078A:q <= 8'h10;
            12'h078B:q <= 8'h1A;
            12'h078C:q <= 8'h18;
            12'h078D:q <= 8'hFF;
            12'h078E:q <= 8'h11;
            12'h078F:q <= 8'h37;
            12'h0790:q <= 8'h48;
            12'h0791:q <= 8'hFF;
            12'h0792:q <= 8'h12;
            12'h0793:q <= 8'h3B;
            12'h0794:q <= 8'h4C;
            12'h0795:q <= 8'hFF;
            12'h0796:q <= 8'h13;
            12'h0797:q <= 8'h52;
            12'h0798:q <= 8'h27;
            12'h0799:q <= 8'hFF;
            12'h079A:q <= 8'h14;
            12'h079B:q <= 8'h58;
            12'h079C:q <= 8'h11;
            12'h079D:q <= 8'hFF;
            12'h079E:q <= 8'h15;
            12'h079F:q <= 8'h3C;
            12'h07A0:q <= 8'h29;
            12'h07A1:q <= 8'hFF;
            12'h07A2:q <= 8'h16;
            12'h07A3:q <= 8'h29;
            12'h07A4:q <= 8'h09;
            12'h07A5:q <= 8'hFF;
            12'h07A6:q <= 8'h17;
            12'h07A7:q <= 8'h2B;
            12'h07A8:q <= 8'h10;
            12'h07A9:q <= 8'hFF;
            12'h07AA:q <= 8'h18;
            12'h07AB:q <= 8'h39;
            12'h07AC:q <= 8'h32;
            12'h07AD:q <= 8'hFF;
            12'h07AE:q <= 8'h19;
            12'h07AF:q <= 8'h3D;
            12'h07B0:q <= 8'h25;
            12'h07B1:q <= 8'hFF;
            12'h07B2:q <= 8'h1A;
            12'h07B3:q <= 8'h53;
            12'h07B4:q <= 8'h49;
            12'h07B5:q <= 8'hFF;
            12'h07B6:q <= 8'h1B;
            12'h07B7:q <= 8'h0F;
            12'h07B8:q <= 8'h0E;
            12'h07B9:q <= 8'hFF;
            12'h07BA:q <= 8'h1C;
            12'h07BB:q <= 8'h20;
            12'h07BC:q <= 8'h50;
            12'h07BD:q <= 8'hFF;
            12'h07BE:q <= 8'h1D;
            12'h07BF:q <= 8'h3E;
            12'h07C0:q <= 8'h2F;
            12'h07C1:q <= 8'hFF;
            12'h07C2:q <= 8'h1E;
            12'h07C3:q <= 8'h0D;
            12'h07C4:q <= 8'h1B;
            12'h07C5:q <= 8'hFF;
            12'h07C6:q <= 8'h1F;
            12'h07C7:q <= 8'h0E;
            12'h07C8:q <= 8'h15;
            12'h07C9:q <= 8'hFF;
            12'h07CA:q <= 8'h20;
            12'h07CB:q <= 8'h03;
            12'h07CC:q <= 8'h35;
            12'h07CD:q <= 8'hFF;
            12'h07CE:q <= 8'h21;
            12'h07CF:q <= 8'h54;
            12'h07D0:q <= 8'h4B;
            12'h07D1:q <= 8'hFF;
            12'h07D2:q <= 8'h22;
            12'h07D3:q <= 8'h28;
            12'h07D4:q <= 8'h3D;
            12'h07D5:q <= 8'hFF;
            12'h07D6:q <= 8'h23;
            12'h07D7:q <= 8'h2E;
            12'h07D8:q <= 8'h16;
            12'h07D9:q <= 8'hFF;
            12'h07DA:q <= 8'h24;
            12'h07DB:q <= 8'h41;
            12'h07DC:q <= 8'h51;
            12'h07DD:q <= 8'hFF;
            12'h07DE:q <= 8'h25;
            12'h07DF:q <= 8'h10;
            12'h07E0:q <= 8'h34;
            12'h07E1:q <= 8'hFF;
            12'h07E2:q <= 8'h26;
            12'h07E3:q <= 8'h00;
            12'h07E4:q <= 8'h14;
            12'h07E5:q <= 8'hFF;
            12'h07E6:q <= 8'h27;
            12'h07E7:q <= 8'h4A;
            12'h07E8:q <= 8'h28;
            12'h07E9:q <= 8'hFF;
            12'h07EA:q <= 8'h28;
            12'h07EB:q <= 8'h51;
            12'h07EC:q <= 8'h06;
            12'h07ED:q <= 8'hFF;
            12'h07EE:q <= 8'h29;
            12'h07EF:q <= 8'h4B;
            12'h07F0:q <= 8'h22;
            12'h07F1:q <= 8'hFF;
            12'h07F2:q <= 8'h2A;
            12'h07F3:q <= 8'h19;
            12'h07F4:q <= 8'h0C;
            12'h07F5:q <= 8'hFF;
            12'h07F6:q <= 8'h2B;
            12'h07F7:q <= 8'h09;
            12'h07F8:q <= 8'h45;
            12'h07F9:q <= 8'hFF;
            12'h07FA:q <= 8'h2C;
            12'h07FB:q <= 8'h50;
            12'h07FC:q <= 8'h1F;
            12'h07FD:q <= 8'hFF;
            12'h07FE:q <= 8'h2D;
            12'h07FF:q <= 8'h12;
            12'h0800:q <= 8'h42;
            12'h0801:q <= 8'hFF;
            12'h0802:q <= 8'h2E;
            12'h0803:q <= 8'h4F;
            12'h0804:q <= 8'h04;
            12'h0805:q <= 8'hFF;
            12'h0806:q <= 8'h2F;
            12'h0807:q <= 8'h36;
            12'h0808:q <= 8'h1A;
            12'h0809:q <= 8'hFF;
            12'h080A:q <= 8'h30;
            12'h080B:q <= 8'h45;
            12'h080C:q <= 8'h57;
            12'h080D:q <= 8'hFF;
            12'h080E:q <= 8'h31;
            12'h080F:q <= 8'h16;
            12'h0810:q <= 8'h33;
            12'h0811:q <= 8'hFF;
            12'h0812:q <= 8'h32;
            12'h0813:q <= 8'h2A;
            12'h0814:q <= 8'h1E;
            12'h0815:q <= 8'hFF;
            12'h0816:q <= 8'h33;
            12'h0817:q <= 8'h34;
            12'h0818:q <= 8'h08;
            12'h0819:q <= 8'hFF;
            12'h081A:q <= 8'h34;
            12'h081B:q <= 8'h22;
            12'h081C:q <= 8'h37;
            12'h081D:q <= 8'hFF;
            12'h081E:q <= 8'h35;
            12'h081F:q <= 8'h07;
            12'h0820:q <= 8'h2B;
            12'h0821:q <= 8'hFF;
            12'h0822:q <= 8'h14;
            12'h0823:q <= 8'h0C;
            12'h0824:q <= 8'h0B;
            12'h0825:q <= 8'h04;
            12'h0826:q <= 8'h0B;
            12'h0827:q <= 8'h0C;
            12'h0828:q <= 8'h14;
            12'h0829:q <= 8'h08;
            12'h082A:q <= 8'hFF;
            12'h082B:q <= 8'h15;
            12'h082C:q <= 8'h12;
            12'h082D:q <= 8'h17;
            12'h082E:q <= 8'h16;
            12'h082F:q <= 8'h17;
            12'h0830:q <= 8'h0E;
            12'h0831:q <= 8'h03;
            12'h0832:q <= 8'h01;
            12'h0833:q <= 8'hFF;
            12'h0834:q <= 8'h16;
            12'h0835:q <= 8'h01;
            12'h0836:q <= 8'h01;
            12'h0837:q <= 8'h13;
            12'h0838:q <= 8'h12;
            12'h0839:q <= 8'h0D;
            12'h083A:q <= 8'h0F;
            12'h083B:q <= 8'h07;
            12'h083C:q <= 8'hFF;
            12'h083D:q <= 8'h17;
            12'h083E:q <= 8'h02;
            12'h083F:q <= 8'h14;
            12'h0840:q <= 8'h02;
            12'h0841:q <= 8'h18;
            12'h0842:q <= 8'h10;
            12'h0843:q <= 8'h11;
            12'h0844:q <= 8'h18;
            12'h0845:q <= 8'hFF;
            12'h0846:q <= 8'h18;
            12'h0847:q <= 8'h0F;
            12'h0848:q <= 8'h03;
            12'h0849:q <= 8'h0D;
            12'h084A:q <= 8'h11;
            12'h084B:q <= 8'h16;
            12'h084C:q <= 8'h0A;
            12'h084D:q <= 8'h02;
            12'h084E:q <= 8'hFF;
            12'h084F:q <= 8'h00;
            12'h0850:q <= 8'h15;
            12'h0851:q <= 8'h09;
            12'h0852:q <= 8'hFF;
            12'h0853:q <= 8'h01;
            12'h0854:q <= 8'h05;
            12'h0855:q <= 8'h10;
            12'h0856:q <= 8'hFF;
            12'h0857:q <= 8'h02;
            12'h0858:q <= 8'h13;
            12'h0859:q <= 8'h0C;
            12'h085A:q <= 8'hFF;
            12'h085B:q <= 8'h03;
            12'h085C:q <= 8'h0E;
            12'h085D:q <= 8'h08;
            12'h085E:q <= 8'hFF;
            12'h085F:q <= 8'h04;
            12'h0860:q <= 8'h00;
            12'h0861:q <= 8'h16;
            12'h0862:q <= 8'hFF;
            12'h0863:q <= 8'h05;
            12'h0864:q <= 8'h18;
            12'h0865:q <= 8'h0F;
            12'h0866:q <= 8'hFF;
            12'h0867:q <= 8'h06;
            12'h0868:q <= 8'h11;
            12'h0869:q <= 8'h18;
            12'h086A:q <= 8'hFF;
            12'h086B:q <= 8'h07;
            12'h086C:q <= 8'h14;
            12'h086D:q <= 8'h11;
            12'h086E:q <= 8'hFF;
            12'h086F:q <= 8'h08;
            12'h0870:q <= 8'h06;
            12'h0871:q <= 8'h05;
            12'h0872:q <= 8'hFF;
            12'h0873:q <= 8'h09;
            12'h0874:q <= 8'h08;
            12'h0875:q <= 8'h02;
            12'h0876:q <= 8'hFF;
            12'h0877:q <= 8'h0A;
            12'h0878:q <= 8'h09;
            12'h0879:q <= 8'h12;
            12'h087A:q <= 8'hFF;
            12'h087B:q <= 8'h0B;
            12'h087C:q <= 8'h0A;
            12'h087D:q <= 8'h15;
            12'h087E:q <= 8'hFF;
            12'h087F:q <= 8'h0C;
            12'h0880:q <= 8'h03;
            12'h0881:q <= 8'h0E;
            12'h0882:q <= 8'hFF;
            12'h0883:q <= 8'h0D;
            12'h0884:q <= 8'h0D;
            12'h0885:q <= 8'h07;
            12'h0886:q <= 8'hFF;
            12'h0887:q <= 8'h0E;
            12'h0888:q <= 8'h0B;
            12'h0889:q <= 8'h00;
            12'h088A:q <= 8'hFF;
            12'h088B:q <= 8'h1E;
            12'h088C:q <= 8'h3A;
            12'h088D:q <= 8'h22;
            12'h088E:q <= 8'h35;
            12'h088F:q <= 8'h01;
            12'h0890:q <= 8'h2A;
            12'h0891:q <= 8'h1A;
            12'h0892:q <= 8'h1B;
            12'h0893:q <= 8'h09;
            12'h0894:q <= 8'h00;
            12'h0895:q <= 8'h3E;
            12'h0896:q <= 8'h23;
            12'h0897:q <= 8'hFF;
            12'h0898:q <= 8'h1F;
            12'h0899:q <= 8'h12;
            12'h089A:q <= 8'h17;
            12'h089B:q <= 8'h24;
            12'h089C:q <= 8'h19;
            12'h089D:q <= 8'h18;
            12'h089E:q <= 8'h0A;
            12'h089F:q <= 8'h25;
            12'h08A0:q <= 8'h3F;
            12'h08A1:q <= 8'h19;
            12'h08A2:q <= 8'h33;
            12'h08A3:q <= 8'h37;
            12'h08A4:q <= 8'hFF;
            12'h08A5:q <= 8'h21;
            12'h08A6:q <= 8'h1D;
            12'h08A7:q <= 8'h02;
            12'h08A8:q <= 8'h3C;
            12'h08A9:q <= 8'h1C;
            12'h08AA:q <= 8'h15;
            12'h08AB:q <= 8'h14;
            12'h08AC:q <= 8'h11;
            12'h08AD:q <= 8'h13;
            12'h08AE:q <= 8'h2A;
            12'h08AF:q <= 8'h39;
            12'h08B0:q <= 8'h2D;
            12'h08B1:q <= 8'hFF;
            12'h08B2:q <= 8'h15;
            12'h08B3:q <= 8'h31;
            12'h08B4:q <= 8'h23;
            12'h08B5:q <= 8'h3D;
            12'h08B6:q <= 8'h21;
            12'h08B7:q <= 8'h23;
            12'h08B8:q <= 8'h08;
            12'h08B9:q <= 8'h0D;
            12'h08BA:q <= 8'h3B;
            12'h08BB:q <= 8'h22;
            12'h08BC:q <= 8'h0D;
            12'h08BD:q <= 8'h16;
            12'h08BE:q <= 8'hFF;
            12'h08BF:q <= 8'h29;
            12'h08C0:q <= 8'h0F;
            12'h08C1:q <= 8'h0B;
            12'h08C2:q <= 8'h3B;
            12'h08C3:q <= 8'h12;
            12'h08C4:q <= 8'h1F;
            12'h08C5:q <= 8'h3F;
            12'h08C6:q <= 8'h2B;
            12'h08C7:q <= 8'h15;
            12'h08C8:q <= 8'h30;
            12'h08C9:q <= 8'h24;
            12'h08CA:q <= 8'h44;
            12'h08CB:q <= 8'hFF;
            12'h08CC:q <= 8'h0C;
            12'h08CD:q <= 8'h44;
            12'h08CE:q <= 8'h3D;
            12'h08CF:q <= 8'h42;
            12'h08D0:q <= 8'h13;
            12'h08D1:q <= 8'h24;
            12'h08D2:q <= 8'h32;
            12'h08D3:q <= 8'h1D;
            12'h08D4:q <= 8'h3A;
            12'h08D5:q <= 8'h25;
            12'h08D6:q <= 8'h11;
            12'h08D7:q <= 8'h3B;
            12'h08D8:q <= 8'hFF;
            12'h08D9:q <= 8'h02;
            12'h08DA:q <= 8'h3C;
            12'h08DB:q <= 8'h20;
            12'h08DC:q <= 8'h18;
            12'h08DD:q <= 8'h15;
            12'h08DE:q <= 8'h43;
            12'h08DF:q <= 8'h06;
            12'h08E0:q <= 8'h43;
            12'h08E1:q <= 8'h44;
            12'h08E2:q <= 8'h40;
            12'h08E3:q <= 8'h1B;
            12'h08E4:q <= 8'h22;
            12'h08E5:q <= 8'hFF;
            12'h08E6:q <= 8'h09;
            12'h08E7:q <= 8'h0E;
            12'h08E8:q <= 8'h34;
            12'h08E9:q <= 8'h20;
            12'h08EA:q <= 8'h0D;
            12'h08EB:q <= 8'h41;
            12'h08EC:q <= 8'h04;
            12'h08ED:q <= 8'h01;
            12'h08EE:q <= 8'h35;
            12'h08EF:q <= 8'h2F;
            12'h08F0:q <= 8'h13;
            12'h08F1:q <= 8'h32;
            12'h08F2:q <= 8'hFF;
            12'h08F3:q <= 8'h2C;
            12'h08F4:q <= 8'h2E;
            12'h08F5:q <= 8'h08;
            12'h08F6:q <= 8'h1E;
            12'h08F7:q <= 8'h08;
            12'h08F8:q <= 8'h21;
            12'h08F9:q <= 8'h2C;
            12'h08FA:q <= 8'h40;
            12'h08FB:q <= 8'h02;
            12'h08FC:q <= 8'h08;
            12'h08FD:q <= 8'h1E;
            12'h08FE:q <= 8'h2E;
            12'h08FF:q <= 8'hFF;
            12'h0900:q <= 8'h35;
            12'h0901:q <= 8'h35;
            12'h0902:q <= 8'h39;
            12'h0903:q <= 8'h29;
            12'h0904:q <= 8'h0B;
            12'h0905:q <= 8'h01;
            12'h0906:q <= 8'h13;
            12'h0907:q <= 8'h2D;
            12'h0908:q <= 8'h26;
            12'h0909:q <= 8'h10;
            12'h090A:q <= 8'h17;
            12'h090B:q <= 8'h31;
            12'h090C:q <= 8'hFF;
            12'h090D:q <= 8'h2A;
            12'h090E:q <= 8'h1C;
            12'h090F:q <= 8'h14;
            12'h0910:q <= 8'h1B;
            12'h0911:q <= 8'h1F;
            12'h0912:q <= 8'h1C;
            12'h0913:q <= 8'h40;
            12'h0914:q <= 8'h06;
            12'h0915:q <= 8'h07;
            12'h0916:q <= 8'h43;
            12'h0917:q <= 8'h1D;
            12'h0918:q <= 8'h47;
            12'h0919:q <= 8'hFF;
            12'h091A:q <= 8'h0B;
            12'h091B:q <= 8'h0C;
            12'h091C:q <= 8'h01;
            12'h091D:q <= 8'h1D;
            12'h091E:q <= 8'h14;
            12'h091F:q <= 8'h19;
            12'h0920:q <= 8'h0B;
            12'h0921:q <= 8'h45;
            12'h0922:q <= 8'h28;
            12'h0923:q <= 8'h26;
            12'h0924:q <= 8'h09;
            12'h0925:q <= 8'h04;
            12'h0926:q <= 8'hFF;
            12'h0927:q <= 8'h26;
            12'h0928:q <= 8'h3B;
            12'h0929:q <= 8'h30;
            12'h092A:q <= 8'h06;
            12'h092B:q <= 8'h2C;
            12'h092C:q <= 8'h3E;
            12'h092D:q <= 8'h33;
            12'h092E:q <= 8'h39;
            12'h092F:q <= 8'h37;
            12'h0930:q <= 8'h2B;
            12'h0931:q <= 8'h03;
            12'h0932:q <= 8'h45;
            12'h0933:q <= 8'hFF;
            12'h0934:q <= 8'h24;
            12'h0935:q <= 8'h46;
            12'h0936:q <= 8'h1E;
            12'h0937:q <= 8'h0E;
            12'h0938:q <= 8'h2F;
            12'h0939:q <= 8'h10;
            12'h093A:q <= 8'h0C;
            12'h093B:q <= 8'h23;
            12'h093C:q <= 8'h31;
            12'h093D:q <= 8'h0A;
            12'h093E:q <= 8'h35;
            12'h093F:q <= 8'h30;
            12'h0940:q <= 8'hFF;
            12'h0941:q <= 8'h12;
            12'h0942:q <= 8'h21;
            12'h0943:q <= 8'h04;
            12'h0944:q <= 8'h41;
            12'h0945:q <= 8'h02;
            12'h0946:q <= 8'h3D;
            12'h0947:q <= 8'h44;
            12'h0948:q <= 8'h1A;
            12'h0949:q <= 8'h32;
            12'h094A:q <= 8'h34;
            12'h094B:q <= 8'h12;
            12'h094C:q <= 8'h33;
            12'h094D:q <= 8'hFF;
            12'h094E:q <= 8'h0F;
            12'h094F:q <= 8'h27;
            12'h0950:q <= 8'h2C;
            12'h0951:q <= 8'h38;
            12'h0952:q <= 8'h00;
            12'h0953:q <= 8'h0D;
            12'h0954:q <= 8'h47;
            12'h0955:q <= 8'h0E;
            12'h0956:q <= 8'h0B;
            12'h0957:q <= 8'h15;
            12'h0958:q <= 8'h28;
            12'h0959:q <= 8'h10;
            12'h095A:q <= 8'hFF;
            12'h095B:q <= 8'h1A;
            12'h095C:q <= 8'h36;
            12'h095D:q <= 8'h1B;
            12'h095E:q <= 8'h39;
            12'h095F:q <= 8'h25;
            12'h0960:q <= 8'h3B;
            12'h0961:q <= 8'h38;
            12'h0962:q <= 8'h21;
            12'h0963:q <= 8'h36;
            12'h0964:q <= 8'h0B;
            12'h0965:q <= 8'h46;
            12'h0966:q <= 8'h36;
            12'h0967:q <= 8'hFF;
            12'h0968:q <= 8'h03;
            12'h0969:q <= 8'h1A;
            12'h096A:q <= 8'h16;
            12'h096B:q <= 8'h44;
            12'h096C:q <= 8'h0A;
            12'h096D:q <= 8'h03;
            12'h096E:q <= 8'h0E;
            12'h096F:q <= 8'h41;
            12'h0970:q <= 8'h19;
            12'h0971:q <= 8'h36;
            12'h0972:q <= 8'h06;
            12'h0973:q <= 8'h25;
            12'h0974:q <= 8'hFF;
            12'h0975:q <= 8'h38;
            12'h0976:q <= 8'h15;
            12'h0977:q <= 8'h07;
            12'h0978:q <= 8'h45;
            12'h0979:q <= 8'h37;
            12'h097A:q <= 8'h2B;
            12'h097B:q <= 8'h2D;
            12'h097C:q <= 8'h04;
            12'h097D:q <= 8'h38;
            12'h097E:q <= 8'h04;
            12'h097F:q <= 8'h1C;
            12'h0980:q <= 8'h3D;
            12'h0981:q <= 8'hFF;
            12'h0982:q <= 8'h39;
            12'h0983:q <= 8'h25;
            12'h0984:q <= 8'h10;
            12'h0985:q <= 8'h46;
            12'h0986:q <= 8'h17;
            12'h0987:q <= 8'h36;
            12'h0988:q <= 8'h45;
            12'h0989:q <= 8'h42;
            12'h098A:q <= 8'h22;
            12'h098B:q <= 8'h3B;
            12'h098C:q <= 8'h47;
            12'h098D:q <= 8'h14;
            12'h098E:q <= 8'hFF;
            12'h098F:q <= 8'h27;
            12'h0990:q <= 8'h06;
            12'h0991:q <= 8'h28;
            12'h0992:q <= 8'h32;
            12'h0993:q <= 8'h28;
            12'h0994:q <= 8'h31;
            12'h0995:q <= 8'h12;
            12'h0996:q <= 8'h27;
            12'h0997:q <= 8'h2C;
            12'h0998:q <= 8'h3D;
            12'h0999:q <= 8'h18;
            12'h099A:q <= 8'h42;
            12'h099B:q <= 8'hFF;
            12'h099C:q <= 8'h20;
            12'h099D:q <= 8'h47;
            12'h099E:q <= 8'h2F;
            12'h099F:q <= 8'h47;
            12'h09A0:q <= 8'h34;
            12'h09A1:q <= 8'h34;
            12'h09A2:q <= 8'h30;
            12'h09A3:q <= 8'h30;
            12'h09A4:q <= 8'h3D;
            12'h09A5:q <= 8'h16;
            12'h09A6:q <= 8'h42;
            12'h09A7:q <= 8'h18;
            12'h09A8:q <= 8'hFF;
            12'h09A9:q <= 8'h3F;
            12'h09AA:q <= 8'h2A;
            12'h09AB:q <= 8'h38;
            12'h09AC:q <= 8'h09;
            12'h09AD:q <= 8'h03;
            12'h09AE:q <= 8'h00;
            12'h09AF:q <= 8'h27;
            12'h09B0:q <= 8'h20;
            12'h09B1:q <= 8'h1E;
            12'h09B2:q <= 8'h05;
            12'h09B3:q <= 8'h38;
            12'h09B4:q <= 8'h08;
            12'h09B5:q <= 8'hFF;
            12'h09B6:q <= 8'h11;
            12'h09B7:q <= 8'h40;
            12'h09B8:q <= 8'h0A;
            12'h09B9:q <= 8'h33;
            12'h09BA:q <= 8'h22;
            12'h09BB:q <= 8'h22;
            12'h09BC:q <= 8'h20;
            12'h09BD:q <= 8'h14;
            12'h09BE:q <= 8'h12;
            12'h09BF:q <= 8'h31;
            12'h09C0:q <= 8'h0F;
            12'h09C1:q <= 8'h34;
            12'h09C2:q <= 8'hFF;
            12'h09C3:q <= 8'h2B;
            12'h09C4:q <= 8'h00;
            12'h09C5:q <= 8'h42;
            12'h09C6:q <= 8'h2E;
            12'h09C7:q <= 8'h23;
            12'h09C8:q <= 8'h25;
            12'h09C9:q <= 8'h46;
            12'h09CA:q <= 8'h24;
            12'h09CB:q <= 8'h0A;
            12'h09CC:q <= 8'h01;
            12'h09CD:q <= 8'h2E;
            12'h09CE:q <= 8'h05;
            12'h09CF:q <= 8'hFF;
            12'h09D0:q <= 8'h06;
            12'h09D1:q <= 8'h19;
            12'h09D2:q <= 8'h05;
            12'h09D3:q <= 8'h26;
            12'h09D4:q <= 8'h04;
            12'h09D5:q <= 8'h3A;
            12'h09D6:q <= 8'h29;
            12'h09D7:q <= 8'h0C;
            12'h09D8:q <= 8'h3C;
            12'h09D9:q <= 8'h29;
            12'h09DA:q <= 8'h07;
            12'h09DB:q <= 8'h28;
            12'h09DC:q <= 8'hFF;
            12'h09DD:q <= 8'h2F;
            12'h09DE:q <= 8'h24;
            12'h09DF:q <= 8'h1F;
            12'h09E0:q <= 8'h16;
            12'h09E1:q <= 8'h11;
            12'h09E2:q <= 8'h28;
            12'h09E3:q <= 8'h16;
            12'h09E4:q <= 8'h2F;
            12'h09E5:q <= 8'h03;
            12'h09E6:q <= 8'h2C;
            12'h09E7:q <= 8'h44;
            12'h09E8:q <= 8'h41;
            12'h09E9:q <= 8'hFF;
            12'h09EA:q <= 8'h17;
            12'h09EB:q <= 8'h13;
            12'h09EC:q <= 8'h03;
            12'h09ED:q <= 8'h0F;
            12'h09EE:q <= 8'h30;
            12'h09EF:q <= 8'h07;
            12'h09F0:q <= 8'h17;
            12'h09F1:q <= 8'h10;
            12'h09F2:q <= 8'h17;
            12'h09F3:q <= 8'h37;
            12'h09F4:q <= 8'h23;
            12'h09F5:q <= 8'h1D;
            12'h09F6:q <= 8'hFF;
            12'h09F7:q <= 8'h43;
            12'h09F8:q <= 8'h3F;
            12'h09F9:q <= 8'h45;
            12'h09FA:q <= 8'h31;
            12'h09FB:q <= 8'h3A;
            12'h09FC:q <= 8'h35;
            12'h09FD:q <= 8'h3C;
            12'h09FE:q <= 8'h46;
            12'h09FF:q <= 8'h05;
            12'h0A00:q <= 8'h0E;
            12'h0A01:q <= 8'h1A;
            12'h0A02:q <= 8'h46;
            12'h0A03:q <= 8'hFF;
            12'h0A04:q <= 8'h3E;
            12'h0A05:q <= 8'h37;
            12'h0A06:q <= 8'h11;
            12'h0A07:q <= 8'h10;
            12'h0A08:q <= 8'h05;
            12'h0A09:q <= 8'h1E;
            12'h0A0A:q <= 8'h42;
            12'h0A0B:q <= 8'h2A;
            12'h0A0C:q <= 8'h16;
            12'h0A0D:q <= 8'h32;
            12'h0A0E:q <= 8'h27;
            12'h0A0F:q <= 8'h0E;
            12'h0A10:q <= 8'hFF;
            12'h0A11:q <= 8'h07;
            12'h0A12:q <= 8'h18;
            12'h0A13:q <= 8'h2D;
            12'h0A14:q <= 8'h3E;
            12'h0A15:q <= 8'h27;
            12'h0A16:q <= 8'h09;
            12'h0A17:q <= 8'h1D;
            12'h0A18:q <= 8'h1C;
            12'h0A19:q <= 8'h29;
            12'h0A1A:q <= 8'h2D;
            12'h0A1B:q <= 8'h21;
            12'h0A1C:q <= 8'h0A;
            12'h0A1D:q <= 8'hFF;
            12'h0A1E:q <= 8'h3A;
            12'h0A1F:q <= 8'h09;
            12'h0A20:q <= 8'h0D;
            12'h0A21:q <= 8'h2A;
            12'h0A22:q <= 8'h07;
            12'h0A23:q <= 8'h05;
            12'h0A24:q <= 8'h37;
            12'h0A25:q <= 8'h47;
            12'h0A26:q <= 8'h0F;
            12'h0A27:q <= 8'h3F;
            12'h0A28:q <= 8'h41;
            12'h0A29:q <= 8'h13;
            12'h0A2A:q <= 8'hFF;
            12'h0A2B:q <= 8'h19;
            12'h0A2C:q <= 8'h3E;
            12'h0A2D:q <= 8'h32;
            12'h0A2E:q <= 8'h3F;
            12'h0A2F:q <= 8'h36;
            12'h0A30:q <= 8'h0F;
            12'h0A31:q <= 8'h1B;
            12'h0A32:q <= 8'h1F;
            12'h0A33:q <= 8'h00;
            12'h0A34:q <= 8'h14;
            12'h0A35:q <= 8'h20;
            12'h0A36:q <= 8'h1C;
            12'h0A37:q <= 8'hFF;
            12'h0A38:q <= 8'h00;
            12'h0A39:q <= 8'h43;
            12'h0A3A:q <= 8'h33;
            12'h0A3B:q <= 8'h2D;
            12'h0A3C:q <= 8'h0C;
            12'h0A3D:q <= 8'h2E;
            12'h0A3E:q <= 8'h02;
            12'h0A3F:q <= 8'h34;
            12'h0A40:q <= 8'h3E;
            12'h0A41:q <= 8'h1F;
            12'h0A42:q <= 8'h3C;
            12'h0A43:q <= 8'h01;
            12'h0A44:q <= 8'hFF;
            12'h0A45:q <= 8'h40;
            12'h0A46:q <= 8'h2B;
            12'h0A47:q <= 8'h29;
            12'h0A48:q <= 8'h2B;
            12'h0A49:q <= 8'h43;
            12'h0A4A:q <= 8'h26;
            12'h0A4B:q <= 8'h39;
            12'h0A4C:q <= 8'h2E;
            12'h0A4D:q <= 8'h33;
            12'h0A4E:q <= 8'h3A;
            12'h0A4F:q <= 8'h02;
            12'h0A50:q <= 8'h0D;
            12'h0A51:q <= 8'hFF;
            12'h0A52:q <= 8'h1B;
            12'h0A53:q <= 8'h41;
            12'h0A54:q <= 8'h26;
            12'h0A55:q <= 8'h1A;
            12'h0A56:q <= 8'h40;
            12'h0A57:q <= 8'h11;
            12'h0A58:q <= 8'h2F;
            12'h0A59:q <= 8'h08;
            12'h0A5A:q <= 8'h18;
            12'h0A5B:q <= 8'h0C;
            12'h0A5C:q <= 8'h45;
            12'h0A5D:q <= 8'h3C;
            12'h0A5E:q <= 8'hFF;
            12'h0A5F:q <= 8'h00;
            12'h0A60:q <= 8'h23;
            12'h0A61:q <= 8'h0D;
            12'h0A62:q <= 8'hFF;
            12'h0A63:q <= 8'h01;
            12'h0A64:q <= 8'h3E;
            12'h0A65:q <= 8'h32;
            12'h0A66:q <= 8'hFF;
            12'h0A67:q <= 8'h02;
            12'h0A68:q <= 8'h08;
            12'h0A69:q <= 8'h21;
            12'h0A6A:q <= 8'hFF;
            12'h0A6B:q <= 8'h03;
            12'h0A6C:q <= 8'h3B;
            12'h0A6D:q <= 8'h34;
            12'h0A6E:q <= 8'hFF;
            12'h0A6F:q <= 8'h04;
            12'h0A70:q <= 8'h00;
            12'h0A71:q <= 8'h2A;
            12'h0A72:q <= 8'hFF;
            12'h0A73:q <= 8'h05;
            12'h0A74:q <= 8'h0C;
            12'h0A75:q <= 8'h10;
            12'h0A76:q <= 8'hFF;
            12'h0A77:q <= 8'h06;
            12'h0A78:q <= 8'h27;
            12'h0A79:q <= 8'h17;
            12'h0A7A:q <= 8'hFF;
            12'h0A7B:q <= 8'h07;
            12'h0A7C:q <= 8'h22;
            12'h0A7D:q <= 8'h1B;
            12'h0A7E:q <= 8'hFF;
            12'h0A7F:q <= 8'h08;
            12'h0A80:q <= 8'h01;
            12'h0A81:q <= 8'h26;
            12'h0A82:q <= 8'hFF;
            12'h0A83:q <= 8'h09;
            12'h0A84:q <= 8'h40;
            12'h0A85:q <= 8'h07;
            12'h0A86:q <= 8'hFF;
            12'h0A87:q <= 8'h0A;
            12'h0A88:q <= 8'h46;
            12'h0A89:q <= 8'h43;
            12'h0A8A:q <= 8'hFF;
            12'h0A8B:q <= 8'h0B;
            12'h0A8C:q <= 8'h1C;
            12'h0A8D:q <= 8'h24;
            12'h0A8E:q <= 8'hFF;
            12'h0A8F:q <= 8'h0C;
            12'h0A90:q <= 8'h45;
            12'h0A91:q <= 8'h05;
            12'h0A92:q <= 8'hFF;
            12'h0A93:q <= 8'h0D;
            12'h0A94:q <= 8'h29;
            12'h0A95:q <= 8'h16;
            12'h0A96:q <= 8'hFF;
            12'h0A97:q <= 8'h0E;
            12'h0A98:q <= 8'h06;
            12'h0A99:q <= 8'h3D;
            12'h0A9A:q <= 8'hFF;
            12'h0A9B:q <= 8'h0F;
            12'h0A9C:q <= 8'h0A;
            12'h0A9D:q <= 8'h19;
            12'h0A9E:q <= 8'hFF;
            12'h0A9F:q <= 8'h10;
            12'h0AA0:q <= 8'h1F;
            12'h0AA1:q <= 8'h1A;
            12'h0AA2:q <= 8'hFF;
            12'h0AA3:q <= 8'h11;
            12'h0AA4:q <= 8'h1E;
            12'h0AA5:q <= 8'h44;
            12'h0AA6:q <= 8'hFF;
            12'h0AA7:q <= 8'h12;
            12'h0AA8:q <= 8'h2F;
            12'h0AA9:q <= 8'h47;
            12'h0AAA:q <= 8'hFF;
            12'h0AAB:q <= 8'h13;
            12'h0AAC:q <= 8'h04;
            12'h0AAD:q <= 8'h2D;
            12'h0AAE:q <= 8'hFF;
            12'h0AAF:q <= 8'h14;
            12'h0AB0:q <= 8'h0B;
            12'h0AB1:q <= 8'h31;
            12'h0AB2:q <= 8'hFF;
            12'h0AB3:q <= 8'h15;
            12'h0AB4:q <= 8'h33;
            12'h0AB5:q <= 8'h03;
            12'h0AB6:q <= 8'hFF;
            12'h0AB7:q <= 8'h16;
            12'h0AB8:q <= 8'h12;
            12'h0AB9:q <= 8'h28;
            12'h0ABA:q <= 8'hFF;
            12'h0ABB:q <= 8'h17;
            12'h0ABC:q <= 8'h1D;
            12'h0ABD:q <= 8'h13;
            12'h0ABE:q <= 8'hFF;
            12'h0ABF:q <= 8'h18;
            12'h0AC0:q <= 8'h0F;
            12'h0AC1:q <= 8'h11;
            12'h0AC2:q <= 8'hFF;
            12'h0AC3:q <= 8'h19;
            12'h0AC4:q <= 8'h39;
            12'h0AC5:q <= 8'h35;
            12'h0AC6:q <= 8'hFF;
            12'h0AC7:q <= 8'h1A;
            12'h0AC8:q <= 8'h15;
            12'h0AC9:q <= 8'h18;
            12'h0ACA:q <= 8'hFF;
            12'h0ACB:q <= 8'h1B;
            12'h0ACC:q <= 8'h37;
            12'h0ACD:q <= 8'h14;
            12'h0ACE:q <= 8'hFF;
            12'h0ACF:q <= 8'h1C;
            12'h0AD0:q <= 8'h02;
            12'h0AD1:q <= 8'h2C;
            12'h0AD2:q <= 8'hFF;
            12'h0AD3:q <= 8'h1D;
            12'h0AD4:q <= 8'h25;
            12'h0AD5:q <= 8'h2E;
            12'h0AD6:q <= 8'hFF;
            12'h0AD7:q <= 8'h1E;
            12'h0AD8:q <= 8'h20;
            12'h0AD9:q <= 8'h3F;
            12'h0ADA:q <= 8'hFF;
            12'h0ADB:q <= 8'h1F;
            12'h0ADC:q <= 8'h3A;
            12'h0ADD:q <= 8'h09;
            12'h0ADE:q <= 8'hFF;
            12'h0ADF:q <= 8'h20;
            12'h0AE0:q <= 8'h36;
            12'h0AE1:q <= 8'h38;
            12'h0AE2:q <= 8'hFF;
            12'h0AE3:q <= 8'h21;
            12'h0AE4:q <= 8'h2B;
            12'h0AE5:q <= 8'h0E;
            12'h0AE6:q <= 8'hFF;
            12'h0AE7:q <= 8'h22;
            12'h0AE8:q <= 8'h41;
            12'h0AE9:q <= 8'h42;
            12'h0AEA:q <= 8'hFF;
            12'h0AEB:q <= 8'h23;
            12'h0AEC:q <= 8'h3C;
            12'h0AED:q <= 8'h30;
            12'h0AEE:q <= 8'hFF;
            12'h0AEF:q <= 8'h24;
            12'h0AF0:q <= 8'h1C;
            12'h0AF1:q <= 8'h30;
            12'h0AF2:q <= 8'hFF;
            12'h0AF3:q <= 8'h25;
            12'h0AF4:q <= 8'h31;
            12'h0AF5:q <= 8'h3F;
            12'h0AF6:q <= 8'hFF;
            12'h0AF7:q <= 8'h26;
            12'h0AF8:q <= 8'h26;
            12'h0AF9:q <= 8'h3B;
            12'h0AFA:q <= 8'hFF;
            12'h0AFB:q <= 8'h27;
            12'h0AFC:q <= 8'h1D;
            12'h0AFD:q <= 8'h15;
            12'h0AFE:q <= 8'hFF;
            12'h0AFF:q <= 8'h28;
            12'h0B00:q <= 8'h19;
            12'h0B01:q <= 8'h1A;
            12'h0B02:q <= 8'hFF;
            12'h0B03:q <= 8'h29;
            12'h0B04:q <= 8'h2E;
            12'h0B05:q <= 8'h09;
            12'h0B06:q <= 8'hFF;
            12'h0B07:q <= 8'h2A;
            12'h0B08:q <= 8'h40;
            12'h0B09:q <= 8'h35;
            12'h0B0A:q <= 8'hFF;
            12'h0B0B:q <= 8'h2B;
            12'h0B0C:q <= 8'h17;
            12'h0B0D:q <= 8'h08;
            12'h0B0E:q <= 8'hFF;
            12'h0B0F:q <= 8'h2C;
            12'h0B10:q <= 8'h0F;
            12'h0B11:q <= 8'h3C;
            12'h0B12:q <= 8'hFF;
            12'h0B13:q <= 8'h2D;
            12'h0B14:q <= 8'h2A;
            12'h0B15:q <= 8'h0D;
            12'h0B16:q <= 8'hFF;
            12'h0B17:q <= 8'h2E;
            12'h0B18:q <= 8'h2C;
            12'h0B19:q <= 8'h0B;
            12'h0B1A:q <= 8'hFF;
            12'h0B1B:q <= 8'h2F;
            12'h0B1C:q <= 8'h21;
            12'h0B1D:q <= 8'h1B;
            12'h0B1E:q <= 8'hFF;
            12'h0B1F:q <= 8'h30;
            12'h0B20:q <= 8'h3E;
            12'h0B21:q <= 8'h33;
            12'h0B22:q <= 8'hFF;
            12'h0B23:q <= 8'h31;
            12'h0B24:q <= 8'h39;
            12'h0B25:q <= 8'h1F;
            12'h0B26:q <= 8'hFF;
            12'h0B27:q <= 8'h32;
            12'h0B28:q <= 8'h27;
            12'h0B29:q <= 8'h18;
            12'h0B2A:q <= 8'hFF;
            12'h0B2B:q <= 8'h33;
            12'h0B2C:q <= 8'h34;
            12'h0B2D:q <= 8'h42;
            12'h0B2E:q <= 8'hFF;
            12'h0B2F:q <= 8'h34;
            12'h0B30:q <= 8'h2B;
            12'h0B31:q <= 8'h20;
            12'h0B32:q <= 8'hFF;
            12'h0B33:q <= 8'h35;
            12'h0B34:q <= 8'h0E;
            12'h0B35:q <= 8'h43;
            12'h0B36:q <= 8'hFF;
            12'h0B37:q <= 8'h36;
            12'h0B38:q <= 8'h11;
            12'h0B39:q <= 8'h46;
            12'h0B3A:q <= 8'hFF;
            12'h0B3B:q <= 8'h37;
            12'h0B3C:q <= 8'h13;
            12'h0B3D:q <= 8'h2F;
            12'h0B3E:q <= 8'hFF;
            12'h0B3F:q <= 8'h38;
            12'h0B40:q <= 8'h02;
            12'h0B41:q <= 8'h14;
            12'h0B42:q <= 8'hFF;
            12'h0B43:q <= 8'h39;
            12'h0B44:q <= 8'h29;
            12'h0B45:q <= 8'h45;
            12'h0B46:q <= 8'hFF;
            12'h0B47:q <= 8'h3A;
            12'h0B48:q <= 8'h05;
            12'h0B49:q <= 8'h0C;
            12'h0B4A:q <= 8'hFF;
            12'h0B4B:q <= 8'h3B;
            12'h0B4C:q <= 8'h3A;
            12'h0B4D:q <= 8'h44;
            12'h0B4E:q <= 8'hFF;
            12'h0B4F:q <= 8'h3C;
            12'h0B50:q <= 8'h04;
            12'h0B51:q <= 8'h23;
            12'h0B52:q <= 8'hFF;
            12'h0B53:q <= 8'h3D;
            12'h0B54:q <= 8'h07;
            12'h0B55:q <= 8'h01;
            12'h0B56:q <= 8'hFF;
            12'h0B57:q <= 8'h3E;
            12'h0B58:q <= 8'h06;
            12'h0B59:q <= 8'h47;
            12'h0B5A:q <= 8'hFF;
            12'h0B5B:q <= 8'h3F;
            12'h0B5C:q <= 8'h12;
            12'h0B5D:q <= 8'h1E;
            12'h0B5E:q <= 8'hFF;
            12'h0B5F:q <= 8'h40;
            12'h0B60:q <= 8'h22;
            12'h0B61:q <= 8'h3D;
            12'h0B62:q <= 8'hFF;
            12'h0B63:q <= 8'h41;
            12'h0B64:q <= 8'h37;
            12'h0B65:q <= 8'h00;
            12'h0B66:q <= 8'hFF;
            12'h0B67:q <= 8'h42;
            12'h0B68:q <= 8'h16;
            12'h0B69:q <= 8'h10;
            12'h0B6A:q <= 8'hFF;
            12'h0B6B:q <= 8'h43;
            12'h0B6C:q <= 8'h25;
            12'h0B6D:q <= 8'h0A;
            12'h0B6E:q <= 8'hFF;
            12'h0B6F:q <= 8'h44;
            12'h0B70:q <= 8'h03;
            12'h0B71:q <= 8'h28;
            12'h0B72:q <= 8'hFF;
            12'h0B73:q <= 8'h45;
            12'h0B74:q <= 8'h36;
            12'h0B75:q <= 8'h38;
            12'h0B76:q <= 8'hFF;
            12'h0B77:q <= 8'h46;
            12'h0B78:q <= 8'h24;
            12'h0B79:q <= 8'h2D;
            12'h0B7A:q <= 8'hFF;
            12'h0B7B:q <= 8'h47;
            12'h0B7C:q <= 8'h32;
            12'h0B7D:q <= 8'h41;
            12'h0B7E:q <= 8'hFF;
            12'h0B7F:q <= 8'h0B;
            12'h0B80:q <= 8'h07;
            12'h0B81:q <= 8'h00;
            12'h0B82:q <= 8'h0E;
            12'h0B83:q <= 8'h06;
            12'h0B84:q <= 8'h05;
            12'h0B85:q <= 8'h04;
            12'h0B86:q <= 8'h04;
            12'h0B87:q <= 8'h0A;
            12'h0B88:q <= 8'h0E;
            12'h0B89:q <= 8'h08;
            12'h0B8A:q <= 8'h0F;
            12'h0B8B:q <= 8'hFF;
            12'h0B8C:q <= 8'h01;
            12'h0B8D:q <= 8'h0D;
            12'h0B8E:q <= 8'h0C;
            12'h0B8F:q <= 8'h03;
            12'h0B90:q <= 8'h04;
            12'h0B91:q <= 8'h0C;
            12'h0B92:q <= 8'h02;
            12'h0B93:q <= 8'h0F;
            12'h0B94:q <= 8'h0D;
            12'h0B95:q <= 8'h03;
            12'h0B96:q <= 8'h11;
            12'h0B97:q <= 8'h05;
            12'h0B98:q <= 8'hFF;
            12'h0B99:q <= 8'h0C;
            12'h0B9A:q <= 8'h0E;
            12'h0B9B:q <= 8'h11;
            12'h0B9C:q <= 8'h00;
            12'h0B9D:q <= 8'h10;
            12'h0B9E:q <= 8'h0A;
            12'h0B9F:q <= 8'h07;
            12'h0BA0:q <= 8'h03;
            12'h0BA1:q <= 8'h01;
            12'h0BA2:q <= 8'h06;
            12'h0BA3:q <= 8'h02;
            12'h0BA4:q <= 8'h02;
            12'h0BA5:q <= 8'hFF;
            12'h0BA6:q <= 8'h09;
            12'h0BA7:q <= 8'h0B;
            12'h0BA8:q <= 8'h05;
            12'h0BA9:q <= 8'h07;
            12'h0BAA:q <= 8'h0C;
            12'h0BAB:q <= 8'h0E;
            12'h0BAC:q <= 8'h0F;
            12'h0BAD:q <= 8'h05;
            12'h0BAE:q <= 8'h00;
            12'h0BAF:q <= 8'h0B;
            12'h0BB0:q <= 8'h0A;
            12'h0BB1:q <= 8'h10;
            12'h0BB2:q <= 8'hFF;
            12'h0BB3:q <= 8'h07;
            12'h0BB4:q <= 8'h10;
            12'h0BB5:q <= 8'h0A;
            12'h0BB6:q <= 8'h05;
            12'h0BB7:q <= 8'h0B;
            12'h0BB8:q <= 8'h10;
            12'h0BB9:q <= 8'h09;
            12'h0BBA:q <= 8'h0E;
            12'h0BBB:q <= 8'h09;
            12'h0BBC:q <= 8'h01;
            12'h0BBD:q <= 8'h10;
            12'h0BBE:q <= 8'h03;
            12'h0BBF:q <= 8'hFF;
            12'h0BC0:q <= 8'h06;
            12'h0BC1:q <= 8'h03;
            12'h0BC2:q <= 8'h09;
            12'h0BC3:q <= 8'h0A;
            12'h0BC4:q <= 8'h01;
            12'h0BC5:q <= 8'h03;
            12'h0BC6:q <= 8'h06;
            12'h0BC7:q <= 8'h08;
            12'h0BC8:q <= 8'h10;
            12'h0BC9:q <= 8'h09;
            12'h0BCA:q <= 8'h0C;
            12'h0BCB:q <= 8'h0D;
            12'h0BCC:q <= 8'hFF;
            12'h0BCD:q <= 8'h08;
            12'h0BCE:q <= 8'h02;
            12'h0BCF:q <= 8'h08;
            12'h0BD0:q <= 8'h09;
            12'h0BD1:q <= 8'h0F;
            12'h0BD2:q <= 8'h01;
            12'h0BD3:q <= 8'h00;
            12'h0BD4:q <= 8'h07;
            12'h0BD5:q <= 8'h0B;
            12'h0BD6:q <= 8'h07;
            12'h0BD7:q <= 8'h0F;
            12'h0BD8:q <= 8'h11;
            12'h0BD9:q <= 8'hFF;
            12'h0BDA:q <= 8'h0E;
            12'h0BDB:q <= 8'h06;
            12'h0BDC:q <= 8'h0F;
            12'h0BDD:q <= 8'h0D;
            12'h0BDE:q <= 8'h08;
            12'h0BDF:q <= 8'h08;
            12'h0BE0:q <= 8'h0B;
            12'h0BE1:q <= 8'h11;
            12'h0BE2:q <= 8'h0C;
            12'h0BE3:q <= 8'h05;
            12'h0BE4:q <= 8'h0D;
            12'h0BE5:q <= 8'h0A;
            12'h0BE6:q <= 8'hFF;
            12'h0BE7:q <= 8'h00;
            12'h0BE8:q <= 8'h04;
            12'h0BE9:q <= 8'h01;
            12'h0BEA:q <= 8'h02;
            12'h0BEB:q <= 8'h11;
            12'h0BEC:q <= 8'h11;
            12'h0BED:q <= 8'h0D;
            12'h0BEE:q <= 8'h06;
            12'h0BEF:q <= 8'h02;
            12'h0BF0:q <= 8'h04;
            12'h0BF1:q <= 8'h00;
            12'h0BF2:q <= 8'h04;
            12'h0BF3:q <= 8'hFF;
            12'h0BF4:q <= 8'h00;
            12'h0BF5:q <= 8'h01;
            12'h0BF6:q <= 8'h07;
            12'h0BF7:q <= 8'hFF;
            12'h0BF8:q <= 8'h01;
            12'h0BF9:q <= 8'h0C;
            12'h0BFA:q <= 8'h03;
            12'h0BFB:q <= 8'hFF;
            12'h0BFC:q <= 8'h02;
            12'h0BFD:q <= 8'h00;
            12'h0BFE:q <= 8'h11;
            12'h0BFF:q <= 8'hFF;
            12'h0C00:q <= 8'h03;
            12'h0C01:q <= 8'h0B;
            12'h0C02:q <= 8'h0D;
            12'h0C03:q <= 8'hFF;
            12'h0C04:q <= 8'h04;
            12'h0C05:q <= 8'h09;
            12'h0C06:q <= 8'h0E;
            12'h0C07:q <= 8'hFF;
            12'h0C08:q <= 8'h05;
            12'h0C09:q <= 8'h05;
            12'h0C0A:q <= 8'h10;
            12'h0C0B:q <= 8'hFF;
            12'h0C0C:q <= 8'h06;
            12'h0C0D:q <= 8'h06;
            12'h0C0E:q <= 8'h0A;
            12'h0C0F:q <= 8'hFF;
            12'h0C10:q <= 8'h07;
            12'h0C11:q <= 8'h08;
            12'h0C12:q <= 8'h02;
            12'h0C13:q <= 8'hFF;
            12'h0C14:q <= 8'h08;
            12'h0C15:q <= 8'h04;
            12'h0C16:q <= 8'h0F;
            12'h0C17:q <= 8'hFF;
            12'h0C18:q <= 8'h09;
            12'h0C19:q <= 8'h0E;
            12'h0C1A:q <= 8'h00;
            12'h0C1B:q <= 8'hFF;
            12'h0C1C:q <= 8'h0A;
            12'h0C1D:q <= 8'h11;
            12'h0C1E:q <= 8'h07;
            12'h0C1F:q <= 8'hFF;
            12'h0C20:q <= 8'h0B;
            12'h0C21:q <= 8'h0B;
            12'h0C22:q <= 8'h0D;
            12'h0C23:q <= 8'hFF;
            12'h0C24:q <= 8'h0C;
            12'h0C25:q <= 8'h08;
            12'h0C26:q <= 8'h05;
            12'h0C27:q <= 8'hFF;
            12'h0C28:q <= 8'h0D;
            12'h0C29:q <= 8'h0A;
            12'h0C2A:q <= 8'h03;
            12'h0C2B:q <= 8'hFF;
            12'h0C2C:q <= 8'h0E;
            12'h0C2D:q <= 8'h06;
            12'h0C2E:q <= 8'h09;
            12'h0C2F:q <= 8'hFF;
            12'h0C30:q <= 8'h0F;
            12'h0C31:q <= 8'h10;
            12'h0C32:q <= 8'h04;
            12'h0C33:q <= 8'hFF;
            12'h0C34:q <= 8'h10;
            12'h0C35:q <= 8'h0F;
            12'h0C36:q <= 8'h02;
            12'h0C37:q <= 8'hFF;
            12'h0C38:q <= 8'h11;
            12'h0C39:q <= 8'h0C;
            12'h0C3A:q <= 8'h01;
            12'h0C3B:q <= 8'hFF;
            12'h0C3C:q <= 8'h00;
            12'h0C3D:q <= 8'h33;
            12'h0C3E:q <= 8'h17;
            12'h0C3F:q <= 8'h1A;
            12'h0C40:q <= 8'h2E;
            12'h0C41:q <= 8'h19;
            12'h0C42:q <= 8'h06;
            12'h0C43:q <= 8'h07;
            12'h0C44:q <= 8'h00;
            12'h0C45:q <= 8'h0D;
            12'h0C46:q <= 8'h27;
            12'h0C47:q <= 8'h13;
            12'h0C48:q <= 8'h30;
            12'h0C49:q <= 8'hFF;
            12'h0C4A:q <= 8'h01;
            12'h0C4B:q <= 8'h3B;
            12'h0C4C:q <= 8'h21;
            12'h0C4D:q <= 8'h0D;
            12'h0C4E:q <= 8'h2C;
            12'h0C4F:q <= 8'h14;
            12'h0C50:q <= 8'h04;
            12'h0C51:q <= 8'h20;
            12'h0C52:q <= 8'h1B;
            12'h0C53:q <= 8'h28;
            12'h0C54:q <= 8'h07;
            12'h0C55:q <= 8'h19;
            12'h0C56:q <= 8'h03;
            12'h0C57:q <= 8'hFF;
            12'h0C58:q <= 8'h02;
            12'h0C59:q <= 8'h11;
            12'h0C5A:q <= 8'h18;
            12'h0C5B:q <= 8'h29;
            12'h0C5C:q <= 8'h1C;
            12'h0C5D:q <= 8'h0E;
            12'h0C5E:q <= 8'h23;
            12'h0C5F:q <= 8'h38;
            12'h0C60:q <= 8'h32;
            12'h0C61:q <= 8'h04;
            12'h0C62:q <= 8'h25;
            12'h0C63:q <= 8'h0F;
            12'h0C64:q <= 8'h0B;
            12'h0C65:q <= 8'hFF;
            12'h0C66:q <= 8'h03;
            12'h0C67:q <= 8'h25;
            12'h0C68:q <= 8'h03;
            12'h0C69:q <= 8'h0C;
            12'h0C6A:q <= 8'h10;
            12'h0C6B:q <= 8'h16;
            12'h0C6C:q <= 8'h31;
            12'h0C6D:q <= 8'h01;
            12'h0C6E:q <= 8'h24;
            12'h0C6F:q <= 8'h3B;
            12'h0C70:q <= 8'h22;
            12'h0C71:q <= 8'h39;
            12'h0C72:q <= 8'h34;
            12'h0C73:q <= 8'hFF;
            12'h0C74:q <= 8'h04;
            12'h0C75:q <= 8'h1F;
            12'h0C76:q <= 8'h09;
            12'h0C77:q <= 8'h30;
            12'h0C78:q <= 8'h3B;
            12'h0C79:q <= 8'h1B;
            12'h0C7A:q <= 8'h37;
            12'h0C7B:q <= 8'h17;
            12'h0C7C:q <= 8'h3A;
            12'h0C7D:q <= 8'h26;
            12'h0C7E:q <= 8'h0E;
            12'h0C7F:q <= 8'h2C;
            12'h0C80:q <= 8'h1A;
            12'h0C81:q <= 8'hFF;
            12'h0C82:q <= 8'h05;
            12'h0C83:q <= 8'h3A;
            12'h0C84:q <= 8'h20;
            12'h0C85:q <= 8'h24;
            12'h0C86:q <= 8'h09;
            12'h0C87:q <= 8'h12;
            12'h0C88:q <= 8'h1E;
            12'h0C89:q <= 8'h33;
            12'h0C8A:q <= 8'h31;
            12'h0C8B:q <= 8'h14;
            12'h0C8C:q <= 8'h05;
            12'h0C8D:q <= 8'h11;
            12'h0C8E:q <= 8'h2A;
            12'h0C8F:q <= 8'hFF;
            12'h0C90:q <= 8'h06;
            12'h0C91:q <= 8'h06;
            12'h0C92:q <= 8'h33;
            12'h0C93:q <= 8'h03;
            12'h0C94:q <= 8'h11;
            12'h0C95:q <= 8'h0B;
            12'h0C96:q <= 8'h35;
            12'h0C97:q <= 8'h2F;
            12'h0C98:q <= 8'h2D;
            12'h0C99:q <= 8'h2B;
            12'h0C9A:q <= 8'h2F;
            12'h0C9B:q <= 8'h1F;
            12'h0C9C:q <= 8'h0A;
            12'h0C9D:q <= 8'hFF;
            12'h0C9E:q <= 8'h07;
            12'h0C9F:q <= 8'h07;
            12'h0CA0:q <= 8'h1F;
            12'h0CA1:q <= 8'h22;
            12'h0CA2:q <= 8'h28;
            12'h0CA3:q <= 8'h0A;
            12'h0CA4:q <= 8'h05;
            12'h0CA5:q <= 8'h15;
            12'h0CA6:q <= 8'h29;
            12'h0CA7:q <= 8'h01;
            12'h0CA8:q <= 8'h15;
            12'h0CA9:q <= 8'h09;
            12'h0CAA:q <= 8'h20;
            12'h0CAB:q <= 8'hFF;
            12'h0CAC:q <= 8'h08;
            12'h0CAD:q <= 8'h0B;
            12'h0CAE:q <= 8'h3B;
            12'h0CAF:q <= 8'h18;
            12'h0CB0:q <= 8'h3A;
            12'h0CB1:q <= 8'h34;
            12'h0CB2:q <= 8'h02;
            12'h0CB3:q <= 8'h32;
            12'h0CB4:q <= 8'h06;
            12'h0CB5:q <= 8'h37;
            12'h0CB6:q <= 8'h16;
            12'h0CB7:q <= 8'h2E;
            12'h0CB8:q <= 8'h36;
            12'h0CB9:q <= 8'hFF;
            12'h0CBA:q <= 8'h09;
            12'h0CBB:q <= 8'h19;
            12'h0CBC:q <= 8'h05;
            12'h0CBD:q <= 8'h25;
            12'h0CBE:q <= 8'h13;
            12'h0CBF:q <= 8'h26;
            12'h0CC0:q <= 8'h1D;
            12'h0CC1:q <= 8'h2B;
            12'h0CC2:q <= 8'h0C;
            12'h0CC3:q <= 8'h1E;
            12'h0CC4:q <= 8'h12;
            12'h0CC5:q <= 8'h38;
            12'h0CC6:q <= 8'h21;
            12'h0CC7:q <= 8'hFF;
            12'h0CC8:q <= 8'h0A;
            12'h0CC9:q <= 8'h1C;
            12'h0CCA:q <= 8'h31;
            12'h0CCB:q <= 8'h2A;
            12'h0CCC:q <= 8'h2D;
            12'h0CCD:q <= 8'h0F;
            12'h0CCE:q <= 8'h39;
            12'h0CCF:q <= 8'h21;
            12'h0CD0:q <= 8'h10;
            12'h0CD1:q <= 8'h35;
            12'h0CD2:q <= 8'h08;
            12'h0CD3:q <= 8'h1C;
            12'h0CD4:q <= 8'h33;
            12'h0CD5:q <= 8'hFF;
            12'h0CD6:q <= 8'h0B;
            12'h0CD7:q <= 8'h20;
            12'h0CD8:q <= 8'h0D;
            12'h0CD9:q <= 8'h27;
            12'h0CDA:q <= 8'h08;
            12'h0CDB:q <= 8'h1F;
            12'h0CDC:q <= 8'h36;
            12'h0CDD:q <= 8'h00;
            12'h0CDE:q <= 8'h1D;
            12'h0CDF:q <= 8'h17;
            12'h0CE0:q <= 8'h18;
            12'h0CE1:q <= 8'h23;
            12'h0CE2:q <= 8'h02;
            12'h0CE3:q <= 8'hFF;
            12'h0CE4:q <= 8'h0C;
            12'h0CE5:q <= 8'h00;
            12'h0CE6:q <= 8'h01;
            12'h0CE7:q <= 8'hFF;
            12'h0CE8:q <= 8'h0D;
            12'h0CE9:q <= 8'h08;
            12'h0CEA:q <= 8'h2F;
            12'h0CEB:q <= 8'hFF;
            12'h0CEC:q <= 8'h0E;
            12'h0CED:q <= 8'h35;
            12'h0CEE:q <= 8'h07;
            12'h0CEF:q <= 8'hFF;
            12'h0CF0:q <= 8'h0F;
            12'h0CF1:q <= 8'h2E;
            12'h0CF2:q <= 8'h2A;
            12'h0CF3:q <= 8'hFF;
            12'h0CF4:q <= 8'h10;
            12'h0CF5:q <= 8'h03;
            12'h0CF6:q <= 8'h14;
            12'h0CF7:q <= 8'hFF;
            12'h0CF8:q <= 8'h11;
            12'h0CF9:q <= 8'h01;
            12'h0CFA:q <= 8'h36;
            12'h0CFB:q <= 8'hFF;
            12'h0CFC:q <= 8'h12;
            12'h0CFD:q <= 8'h30;
            12'h0CFE:q <= 8'h1E;
            12'h0CFF:q <= 8'hFF;
            12'h0D00:q <= 8'h13;
            12'h0D01:q <= 8'h24;
            12'h0D02:q <= 8'h10;
            12'h0D03:q <= 8'hFF;
            12'h0D04:q <= 8'h14;
            12'h0D05:q <= 8'h37;
            12'h0D06:q <= 8'h25;
            12'h0D07:q <= 8'hFF;
            12'h0D08:q <= 8'h15;
            12'h0D09:q <= 8'h31;
            12'h0D0A:q <= 8'h26;
            12'h0D0B:q <= 8'hFF;
            12'h0D0C:q <= 8'h16;
            12'h0D0D:q <= 8'h28;
            12'h0D0E:q <= 8'h1C;
            12'h0D0F:q <= 8'hFF;
            12'h0D10:q <= 8'h17;
            12'h0D11:q <= 8'h23;
            12'h0D12:q <= 8'h0E;
            12'h0D13:q <= 8'hFF;
            12'h0D14:q <= 8'h18;
            12'h0D15:q <= 8'h29;
            12'h0D16:q <= 8'h32;
            12'h0D17:q <= 8'hFF;
            12'h0D18:q <= 8'h19;
            12'h0D19:q <= 8'h0F;
            12'h0D1A:q <= 8'h2C;
            12'h0D1B:q <= 8'hFF;
            12'h0D1C:q <= 8'h1A;
            12'h0D1D:q <= 8'h21;
            12'h0D1E:q <= 8'h23;
            12'h0D1F:q <= 8'hFF;
            12'h0D20:q <= 8'h1B;
            12'h0D21:q <= 8'h0E;
            12'h0D22:q <= 8'h2B;
            12'h0D23:q <= 8'hFF;
            12'h0D24:q <= 8'h1C;
            12'h0D25:q <= 8'h1D;
            12'h0D26:q <= 8'h15;
            12'h0D27:q <= 8'hFF;
            12'h0D28:q <= 8'h1D;
            12'h0D29:q <= 8'h12;
            12'h0D2A:q <= 8'h27;
            12'h0D2B:q <= 8'hFF;
            12'h0D2C:q <= 8'h1E;
            12'h0D2D:q <= 8'h04;
            12'h0D2E:q <= 8'h1B;
            12'h0D2F:q <= 8'hFF;
            12'h0D30:q <= 8'h1F;
            12'h0D31:q <= 8'h32;
            12'h0D32:q <= 8'h08;
            12'h0D33:q <= 8'hFF;
            12'h0D34:q <= 8'h20;
            12'h0D35:q <= 8'h26;
            12'h0D36:q <= 8'h37;
            12'h0D37:q <= 8'hFF;
            12'h0D38:q <= 8'h21;
            12'h0D39:q <= 8'h2B;
            12'h0D3A:q <= 8'h0B;
            12'h0D3B:q <= 8'hFF;
            12'h0D3C:q <= 8'h22;
            12'h0D3D:q <= 8'h10;
            12'h0D3E:q <= 8'h11;
            12'h0D3F:q <= 8'hFF;
            12'h0D40:q <= 8'h23;
            12'h0D41:q <= 8'h1E;
            12'h0D42:q <= 8'h06;
            12'h0D43:q <= 8'hFF;
            12'h0D44:q <= 8'h24;
            12'h0D45:q <= 8'h15;
            12'h0D46:q <= 8'h2D;
            12'h0D47:q <= 8'hFF;
            12'h0D48:q <= 8'h25;
            12'h0D49:q <= 8'h27;
            12'h0D4A:q <= 8'h19;
            12'h0D4B:q <= 8'hFF;
            12'h0D4C:q <= 8'h26;
            12'h0D4D:q <= 8'h0A;
            12'h0D4E:q <= 8'h12;
            12'h0D4F:q <= 8'hFF;
            12'h0D50:q <= 8'h27;
            12'h0D51:q <= 8'h02;
            12'h0D52:q <= 8'h00;
            12'h0D53:q <= 8'hFF;
            12'h0D54:q <= 8'h28;
            12'h0D55:q <= 8'h0D;
            12'h0D56:q <= 8'h34;
            12'h0D57:q <= 8'hFF;
            12'h0D58:q <= 8'h29;
            12'h0D59:q <= 8'h2D;
            12'h0D5A:q <= 8'h2E;
            12'h0D5B:q <= 8'hFF;
            12'h0D5C:q <= 8'h2A;
            12'h0D5D:q <= 8'h09;
            12'h0D5E:q <= 8'h0A;
            12'h0D5F:q <= 8'hFF;
            12'h0D60:q <= 8'h2B;
            12'h0D61:q <= 8'h39;
            12'h0D62:q <= 8'h35;
            12'h0D63:q <= 8'hFF;
            12'h0D64:q <= 8'h2C;
            12'h0D65:q <= 8'h14;
            12'h0D66:q <= 8'h0C;
            12'h0D67:q <= 8'hFF;
            12'h0D68:q <= 8'h2D;
            12'h0D69:q <= 8'h18;
            12'h0D6A:q <= 8'h30;
            12'h0D6B:q <= 8'hFF;
            12'h0D6C:q <= 8'h2E;
            12'h0D6D:q <= 8'h38;
            12'h0D6E:q <= 8'h29;
            12'h0D6F:q <= 8'hFF;
            12'h0D70:q <= 8'h2F;
            12'h0D71:q <= 8'h13;
            12'h0D72:q <= 8'h02;
            12'h0D73:q <= 8'hFF;
            12'h0D74:q <= 8'h30;
            12'h0D75:q <= 8'h2A;
            12'h0D76:q <= 8'h16;
            12'h0D77:q <= 8'hFF;
            12'h0D78:q <= 8'h31;
            12'h0D79:q <= 8'h36;
            12'h0D7A:q <= 8'h39;
            12'h0D7B:q <= 8'hFF;
            12'h0D7C:q <= 8'h32;
            12'h0D7D:q <= 8'h2F;
            12'h0D7E:q <= 8'h13;
            12'h0D7F:q <= 8'hFF;
            12'h0D80:q <= 8'h33;
            12'h0D81:q <= 8'h34;
            12'h0D82:q <= 8'h24;
            12'h0D83:q <= 8'hFF;
            12'h0D84:q <= 8'h34;
            12'h0D85:q <= 8'h22;
            12'h0D86:q <= 8'h3A;
            12'h0D87:q <= 8'hFF;
            12'h0D88:q <= 8'h35;
            12'h0D89:q <= 8'h17;
            12'h0D8A:q <= 8'h28;
            12'h0D8B:q <= 8'hFF;
            12'h0D8C:q <= 8'h36;
            12'h0D8D:q <= 8'h1A;
            12'h0D8E:q <= 8'h1A;
            12'h0D8F:q <= 8'hFF;
            12'h0D90:q <= 8'h37;
            12'h0D91:q <= 8'h16;
            12'h0D92:q <= 8'h1D;
            12'h0D93:q <= 8'hFF;
            12'h0D94:q <= 8'h38;
            12'h0D95:q <= 8'h0C;
            12'h0D96:q <= 8'h0F;
            12'h0D97:q <= 8'hFF;
            12'h0D98:q <= 8'h39;
            12'h0D99:q <= 8'h05;
            12'h0D9A:q <= 8'h22;
            12'h0D9B:q <= 8'hFF;
            12'h0D9C:q <= 8'h3A;
            12'h0D9D:q <= 8'h1B;
            12'h0D9E:q <= 8'h04;
            12'h0D9F:q <= 8'hFF;
            12'h0DA0:q <= 8'h3B;
            12'h0DA1:q <= 8'h2C;
            12'h0DA2:q <= 8'h38;
            12'h0DA3:q <= 8'hFF;
            12'h0DA4:q <= 8'h00;
            12'h0DA5:q <= 8'h2E;
            12'h0DA6:q <= 8'h2F;
            12'h0DA7:q <= 8'hFF;
            12'h0DA8:q <= 8'h01;
            12'h0DA9:q <= 8'h14;
            12'h0DAA:q <= 8'h2E;
            12'h0DAB:q <= 8'hFF;
            12'h0DAC:q <= 8'h02;
            12'h0DAD:q <= 8'h35;
            12'h0DAE:q <= 8'h05;
            12'h0DAF:q <= 8'hFF;
            12'h0DB0:q <= 8'h03;
            12'h0DB1:q <= 8'h0C;
            12'h0DB2:q <= 8'h39;
            12'h0DB3:q <= 8'hFF;
            12'h0DB4:q <= 8'h04;
            12'h0DB5:q <= 8'h29;
            12'h0DB6:q <= 8'h2A;
            12'h0DB7:q <= 8'hFF;
            12'h0DB8:q <= 8'h05;
            12'h0DB9:q <= 8'h22;
            12'h0DBA:q <= 8'h0D;
            12'h0DBB:q <= 8'hFF;
            12'h0DBC:q <= 8'h06;
            12'h0DBD:q <= 8'h05;
            12'h0DBE:q <= 8'h12;
            12'h0DBF:q <= 8'hFF;
            12'h0DC0:q <= 8'h07;
            12'h0DC1:q <= 8'h13;
            12'h0DC2:q <= 8'h3A;
            12'h0DC3:q <= 8'hFF;
            12'h0DC4:q <= 8'h08;
            12'h0DC5:q <= 8'h18;
            12'h0DC6:q <= 8'h23;
            12'h0DC7:q <= 8'hFF;
            12'h0DC8:q <= 8'h09;
            12'h0DC9:q <= 8'h06;
            12'h0DCA:q <= 8'h22;
            12'h0DCB:q <= 8'hFF;
            12'h0DCC:q <= 8'h0A;
            12'h0DCD:q <= 8'h36;
            12'h0DCE:q <= 8'h16;
            12'h0DCF:q <= 8'hFF;
            12'h0DD0:q <= 8'h0B;
            12'h0DD1:q <= 8'h0F;
            12'h0DD2:q <= 8'h24;
            12'h0DD3:q <= 8'hFF;
            12'h0DD4:q <= 8'h0C;
            12'h0DD5:q <= 8'h04;
            12'h0DD6:q <= 8'h1B;
            12'h0DD7:q <= 8'hFF;
            12'h0DD8:q <= 8'h0D;
            12'h0DD9:q <= 8'h1D;
            12'h0DDA:q <= 8'h20;
            12'h0DDB:q <= 8'hFF;
            12'h0DDC:q <= 8'h0E;
            12'h0DDD:q <= 8'h16;
            12'h0DDE:q <= 8'h33;
            12'h0DDF:q <= 8'hFF;
            12'h0DE0:q <= 8'h0F;
            12'h0DE1:q <= 8'h2A;
            12'h0DE2:q <= 8'h31;
            12'h0DE3:q <= 8'hFF;
            12'h0DE4:q <= 8'h10;
            12'h0DE5:q <= 8'h0D;
            12'h0DE6:q <= 8'h2D;
            12'h0DE7:q <= 8'hFF;
            12'h0DE8:q <= 8'h11;
            12'h0DE9:q <= 8'h0E;
            12'h0DEA:q <= 8'h1A;
            12'h0DEB:q <= 8'hFF;
            12'h0DEC:q <= 8'h12;
            12'h0DED:q <= 8'h11;
            12'h0DEE:q <= 8'h04;
            12'h0DEF:q <= 8'hFF;
            12'h0DF0:q <= 8'h13;
            12'h0DF1:q <= 8'h00;
            12'h0DF2:q <= 8'h00;
            12'h0DF3:q <= 8'hFF;
            12'h0DF4:q <= 8'h14;
            12'h0DF5:q <= 8'h20;
            12'h0DF6:q <= 8'h36;
            12'h0DF7:q <= 8'hFF;
            12'h0DF8:q <= 8'h15;
            12'h0DF9:q <= 8'h1A;
            12'h0DFA:q <= 8'h15;
            12'h0DFB:q <= 8'hFF;
            12'h0DFC:q <= 8'h16;
            12'h0DFD:q <= 8'h0B;
            12'h0DFE:q <= 8'h0E;
            12'h0DFF:q <= 8'hFF;
            12'h0E00:q <= 8'h17;
            12'h0E01:q <= 8'h39;
            12'h0E02:q <= 8'h06;
            12'h0E03:q <= 8'hFF;
            12'h0E04:q <= 8'h18;
            12'h0E05:q <= 8'h2D;
            12'h0E06:q <= 8'h13;
            12'h0E07:q <= 8'hFF;
            12'h0E08:q <= 8'h19;
            12'h0E09:q <= 8'h02;
            12'h0E0A:q <= 8'h0A;
            12'h0E0B:q <= 8'hFF;
            12'h0E0C:q <= 8'h1A;
            12'h0E0D:q <= 8'h10;
            12'h0E0E:q <= 8'h1E;
            12'h0E0F:q <= 8'hFF;
            12'h0E10:q <= 8'h1B;
            12'h0E11:q <= 8'h15;
            12'h0E12:q <= 8'h29;
            12'h0E13:q <= 8'hFF;
            12'h0E14:q <= 8'h1C;
            12'h0E15:q <= 8'h12;
            12'h0E16:q <= 8'h07;
            12'h0E17:q <= 8'hFF;
            12'h0E18:q <= 8'h1D;
            12'h0E19:q <= 8'h3A;
            12'h0E1A:q <= 8'h18;
            12'h0E1B:q <= 8'hFF;
            12'h0E1C:q <= 8'h1E;
            12'h0E1D:q <= 8'h2C;
            12'h0E1E:q <= 8'h14;
            12'h0E1F:q <= 8'hFF;
            12'h0E20:q <= 8'h1F;
            12'h0E21:q <= 8'h24;
            12'h0E22:q <= 8'h1D;
            12'h0E23:q <= 8'hFF;
            12'h0E24:q <= 8'h20;
            12'h0E25:q <= 8'h30;
            12'h0E26:q <= 8'h26;
            12'h0E27:q <= 8'hFF;
            12'h0E28:q <= 8'h21;
            12'h0E29:q <= 8'h27;
            12'h0E2A:q <= 8'h2C;
            12'h0E2B:q <= 8'hFF;
            12'h0E2C:q <= 8'h22;
            12'h0E2D:q <= 8'h0A;
            12'h0E2E:q <= 8'h09;
            12'h0E2F:q <= 8'hFF;
            12'h0E30:q <= 8'h23;
            12'h0E31:q <= 8'h28;
            12'h0E32:q <= 8'h34;
            12'h0E33:q <= 8'hFF;
            12'h0E34:q <= 8'h24;
            12'h0E35:q <= 8'h1B;
            12'h0E36:q <= 8'h2B;
            12'h0E37:q <= 8'hFF;
            12'h0E38:q <= 8'h25;
            12'h0E39:q <= 8'h1E;
            12'h0E3A:q <= 8'h0B;
            12'h0E3B:q <= 8'hFF;
            12'h0E3C:q <= 8'h26;
            12'h0E3D:q <= 8'h25;
            12'h0E3E:q <= 8'h19;
            12'h0E3F:q <= 8'hFF;
            12'h0E40:q <= 8'h27;
            12'h0E41:q <= 8'h07;
            12'h0E42:q <= 8'h25;
            12'h0E43:q <= 8'hFF;
            12'h0E44:q <= 8'h28;
            12'h0E45:q <= 8'h38;
            12'h0E46:q <= 8'h1F;
            12'h0E47:q <= 8'hFF;
            12'h0E48:q <= 8'h29;
            12'h0E49:q <= 8'h34;
            12'h0E4A:q <= 8'h3B;
            12'h0E4B:q <= 8'hFF;
            12'h0E4C:q <= 8'h2A;
            12'h0E4D:q <= 8'h26;
            12'h0E4E:q <= 8'h10;
            12'h0E4F:q <= 8'hFF;
            12'h0E50:q <= 8'h2B;
            12'h0E51:q <= 8'h09;
            12'h0E52:q <= 8'h0C;
            12'h0E53:q <= 8'hFF;
            12'h0E54:q <= 8'h2C;
            12'h0E55:q <= 8'h21;
            12'h0E56:q <= 8'h35;
            12'h0E57:q <= 8'hFF;
            12'h0E58:q <= 8'h2D;
            12'h0E59:q <= 8'h19;
            12'h0E5A:q <= 8'h1C;
            12'h0E5B:q <= 8'hFF;
            12'h0E5C:q <= 8'h2E;
            12'h0E5D:q <= 8'h03;
            12'h0E5E:q <= 8'h37;
            12'h0E5F:q <= 8'hFF;
            12'h0E60:q <= 8'h2F;
            12'h0E61:q <= 8'h08;
            12'h0E62:q <= 8'h0F;
            12'h0E63:q <= 8'hFF;
            12'h0E64:q <= 8'h30;
            12'h0E65:q <= 8'h23;
            12'h0E66:q <= 8'h11;
            12'h0E67:q <= 8'hFF;
            12'h0E68:q <= 8'h31;
            12'h0E69:q <= 8'h2B;
            12'h0E6A:q <= 8'h38;
            12'h0E6B:q <= 8'hFF;
            12'h0E6C:q <= 8'h32;
            12'h0E6D:q <= 8'h3B;
            12'h0E6E:q <= 8'h08;
            12'h0E6F:q <= 8'hFF;
            12'h0E70:q <= 8'h33;
            12'h0E71:q <= 8'h01;
            12'h0E72:q <= 8'h27;
            12'h0E73:q <= 8'hFF;
            12'h0E74:q <= 8'h34;
            12'h0E75:q <= 8'h32;
            12'h0E76:q <= 8'h01;
            12'h0E77:q <= 8'hFF;
            12'h0E78:q <= 8'h35;
            12'h0E79:q <= 8'h1C;
            12'h0E7A:q <= 8'h21;
            12'h0E7B:q <= 8'hFF;
            12'h0E7C:q <= 8'h36;
            12'h0E7D:q <= 8'h2F;
            12'h0E7E:q <= 8'h03;
            12'h0E7F:q <= 8'hFF;
            12'h0E80:q <= 8'h37;
            12'h0E81:q <= 8'h17;
            12'h0E82:q <= 8'h17;
            12'h0E83:q <= 8'hFF;
            12'h0E84:q <= 8'h38;
            12'h0E85:q <= 8'h33;
            12'h0E86:q <= 8'h30;
            12'h0E87:q <= 8'hFF;
            12'h0E88:q <= 8'h39;
            12'h0E89:q <= 8'h1F;
            12'h0E8A:q <= 8'h02;
            12'h0E8B:q <= 8'hFF;
            12'h0E8C:q <= 8'h3A;
            12'h0E8D:q <= 8'h37;
            12'h0E8E:q <= 8'h28;
            12'h0E8F:q <= 8'hFF;
            12'h0E90:q <= 8'h3B;
            12'h0E91:q <= 8'h31;
            12'h0E92:q <= 8'h32;
            12'h0E93:q <= 8'hFF;
            12'h0E94:q <= 8'h00;
            12'h0E95:q <= 8'h0E;
            12'h0E96:q <= 8'h08;
            12'h0E97:q <= 8'h03;
            12'h0E98:q <= 8'h0B;
            12'h0E99:q <= 8'h05;
            12'h0E9A:q <= 8'h01;
            12'h0E9B:q <= 8'h07;
            12'h0E9C:q <= 8'h06;
            12'h0E9D:q <= 8'h09;
            12'h0E9E:q <= 8'h01;
            12'h0E9F:q <= 8'h00;
            12'h0EA0:q <= 8'h0C;
            12'h0EA1:q <= 8'hFF;
            12'h0EA2:q <= 8'h01;
            12'h0EA3:q <= 8'h02;
            12'h0EA4:q <= 8'h01;
            12'h0EA5:q <= 8'h0D;
            12'h0EA6:q <= 8'h00;
            12'h0EA7:q <= 8'h0C;
            12'h0EA8:q <= 8'h02;
            12'h0EA9:q <= 8'h04;
            12'h0EAA:q <= 8'h04;
            12'h0EAB:q <= 8'h0D;
            12'h0EAC:q <= 8'h0B;
            12'h0EAD:q <= 8'h08;
            12'h0EAE:q <= 8'h03;
            12'h0EAF:q <= 8'hFF;
            12'h0EB0:q <= 8'h02;
            12'h0EB1:q <= 8'h04;
            12'h0EB2:q <= 8'h09;
            12'h0EB3:q <= 8'h0E;
            12'h0EB4:q <= 8'h0A;
            12'h0EB5:q <= 8'h09;
            12'h0EB6:q <= 8'h06;
            12'h0EB7:q <= 8'h08;
            12'h0EB8:q <= 8'h02;
            12'h0EB9:q <= 8'h07;
            12'h0EBA:q <= 8'h0E;
            12'h0EBB:q <= 8'h05;
            12'h0EBC:q <= 8'h0A;
            12'h0EBD:q <= 8'hFF;
            12'h0EBE:q <= 8'h03;
            12'h0EBF:q <= 8'h0C;
            12'h0EC0:q <= 8'h04;
            12'h0EC1:q <= 8'hFF;
            12'h0EC2:q <= 8'h04;
            12'h0EC3:q <= 8'h0D;
            12'h0EC4:q <= 8'h02;
            12'h0EC5:q <= 8'hFF;
            12'h0EC6:q <= 8'h05;
            12'h0EC7:q <= 8'h05;
            12'h0EC8:q <= 8'h06;
            12'h0EC9:q <= 8'hFF;
            12'h0ECA:q <= 8'h06;
            12'h0ECB:q <= 8'h09;
            12'h0ECC:q <= 8'h05;
            12'h0ECD:q <= 8'hFF;
            12'h0ECE:q <= 8'h07;
            12'h0ECF:q <= 8'h03;
            12'h0ED0:q <= 8'h0C;
            12'h0ED1:q <= 8'hFF;
            12'h0ED2:q <= 8'h08;
            12'h0ED3:q <= 8'h0B;
            12'h0ED4:q <= 8'h0B;
            12'h0ED5:q <= 8'hFF;
            12'h0ED6:q <= 8'h09;
            12'h0ED7:q <= 8'h07;
            12'h0ED8:q <= 8'h07;
            12'h0ED9:q <= 8'hFF;
            12'h0EDA:q <= 8'h0A;
            12'h0EDB:q <= 8'h01;
            12'h0EDC:q <= 8'h0D;
            12'h0EDD:q <= 8'hFF;
            12'h0EDE:q <= 8'h0B;
            12'h0EDF:q <= 8'h00;
            12'h0EE0:q <= 8'h00;
            12'h0EE1:q <= 8'hFF;
            12'h0EE2:q <= 8'h0C;
            12'h0EE3:q <= 8'h06;
            12'h0EE4:q <= 8'h0A;
            12'h0EE5:q <= 8'hFF;
            12'h0EE6:q <= 8'h0D;
            12'h0EE7:q <= 8'h08;
            12'h0EE8:q <= 8'h0E;
            12'h0EE9:q <= 8'hFF;
            12'h0EEA:q <= 8'h0E;
            12'h0EEB:q <= 8'h0A;
            12'h0EEC:q <= 8'h03;
            12'h0EED:q <= 8'hFF;
            12'h0EEE:q <= 8'h00;
            12'h0EEF:q <= 8'h0D;
            12'h0EF0:q <= 8'h01;
            12'h0EF1:q <= 8'hFF;
            12'h0EF2:q <= 8'h01;
            12'h0EF3:q <= 8'h03;
            12'h0EF4:q <= 8'h0A;
            12'h0EF5:q <= 8'hFF;
            12'h0EF6:q <= 8'h02;
            12'h0EF7:q <= 8'h0C;
            12'h0EF8:q <= 8'h0E;
            12'h0EF9:q <= 8'hFF;
            12'h0EFA:q <= 8'h03;
            12'h0EFB:q <= 8'h08;
            12'h0EFC:q <= 8'h00;
            12'h0EFD:q <= 8'hFF;
            12'h0EFE:q <= 8'h04;
            12'h0EFF:q <= 8'h07;
            12'h0F00:q <= 8'h02;
            12'h0F01:q <= 8'hFF;
            12'h0F02:q <= 8'h05;
            12'h0F03:q <= 8'h0A;
            12'h0F04:q <= 8'h0C;
            12'h0F05:q <= 8'hFF;
            12'h0F06:q <= 8'h06;
            12'h0F07:q <= 8'h02;
            12'h0F08:q <= 8'h0B;
            12'h0F09:q <= 8'hFF;
            12'h0F0A:q <= 8'h07;
            12'h0F0B:q <= 8'h01;
            12'h0F0C:q <= 8'h06;
            12'h0F0D:q <= 8'hFF;
            12'h0F0E:q <= 8'h08;
            12'h0F0F:q <= 8'h00;
            12'h0F10:q <= 8'h07;
            12'h0F11:q <= 8'hFF;
            12'h0F12:q <= 8'h09;
            12'h0F13:q <= 8'h0B;
            12'h0F14:q <= 8'h05;
            12'h0F15:q <= 8'hFF;
            12'h0F16:q <= 8'h0A;
            12'h0F17:q <= 8'h0E;
            12'h0F18:q <= 8'h03;
            12'h0F19:q <= 8'hFF;
            12'h0F1A:q <= 8'h0B;
            12'h0F1B:q <= 8'h09;
            12'h0F1C:q <= 8'h08;
            12'h0F1D:q <= 8'hFF;
            12'h0F1E:q <= 8'h0C;
            12'h0F1F:q <= 8'h05;
            12'h0F20:q <= 8'h0D;
            12'h0F21:q <= 8'hFF;
            12'h0F22:q <= 8'h0D;
            12'h0F23:q <= 8'h06;
            12'h0F24:q <= 8'h04;
            12'h0F25:q <= 8'hFF;
            12'h0F26:q <= 8'h0E;
            12'h0F27:q <= 8'h04;
            12'h0F28:q <= 8'h09;
            12'h0F29:q <= 8'hFF;
            12'h0F2A:q <= 8'h00;
            12'h0F2B:q <= 8'h28;
            12'h0F2C:q <= 8'h1A;
            12'h0F2D:q <= 8'h1F;
            12'h0F2E:q <= 8'h18;
            12'h0F2F:q <= 8'h28;
            12'h0F30:q <= 8'h0C;
            12'h0F31:q <= 8'h17;
            12'h0F32:q <= 8'h1D;
            12'h0F33:q <= 8'h16;
            12'h0F34:q <= 8'h0B;
            12'h0F35:q <= 8'h27;
            12'h0F36:q <= 8'hFF;
            12'h0F37:q <= 8'h01;
            12'h0F38:q <= 8'h13;
            12'h0F39:q <= 8'h2B;
            12'h0F3A:q <= 8'h2A;
            12'h0F3B:q <= 8'h09;
            12'h0F3C:q <= 8'h25;
            12'h0F3D:q <= 8'h2C;
            12'h0F3E:q <= 8'h02;
            12'h0F3F:q <= 8'h0A;
            12'h0F40:q <= 8'h2A;
            12'h0F41:q <= 8'h15;
            12'h0F42:q <= 8'h20;
            12'h0F43:q <= 8'hFF;
            12'h0F44:q <= 8'h02;
            12'h0F45:q <= 8'h20;
            12'h0F46:q <= 8'h0C;
            12'h0F47:q <= 8'h15;
            12'h0F48:q <= 8'h16;
            12'h0F49:q <= 8'h02;
            12'h0F4A:q <= 8'h04;
            12'h0F4B:q <= 8'h11;
            12'h0F4C:q <= 8'h00;
            12'h0F4D:q <= 8'h2B;
            12'h0F4E:q <= 8'h09;
            12'h0F4F:q <= 8'h22;
            12'h0F50:q <= 8'hFF;
            12'h0F51:q <= 8'h03;
            12'h0F52:q <= 8'h1E;
            12'h0F53:q <= 8'h0E;
            12'h0F54:q <= 8'h00;
            12'h0F55:q <= 8'h11;
            12'h0F56:q <= 8'h01;
            12'h0F57:q <= 8'h20;
            12'h0F58:q <= 8'h2A;
            12'h0F59:q <= 8'h10;
            12'h0F5A:q <= 8'h23;
            12'h0F5B:q <= 8'h11;
            12'h0F5C:q <= 8'h24;
            12'h0F5D:q <= 8'hFF;
            12'h0F5E:q <= 8'h04;
            12'h0F5F:q <= 8'h15;
            12'h0F60:q <= 8'h16;
            12'h0F61:q <= 8'h13;
            12'h0F62:q <= 8'h0E;
            12'h0F63:q <= 8'h08;
            12'h0F64:q <= 8'h2B;
            12'h0F65:q <= 8'h09;
            12'h0F66:q <= 8'h0D;
            12'h0F67:q <= 8'h0F;
            12'h0F68:q <= 8'h1F;
            12'h0F69:q <= 8'h0A;
            12'h0F6A:q <= 8'hFF;
            12'h0F6B:q <= 8'h05;
            12'h0F6C:q <= 8'h23;
            12'h0F6D:q <= 8'h1D;
            12'h0F6E:q <= 8'h24;
            12'h0F6F:q <= 8'h29;
            12'h0F70:q <= 8'h05;
            12'h0F71:q <= 8'h05;
            12'h0F72:q <= 8'h03;
            12'h0F73:q <= 8'h0B;
            12'h0F74:q <= 8'h06;
            12'h0F75:q <= 8'h14;
            12'h0F76:q <= 8'h17;
            12'h0F77:q <= 8'hFF;
            12'h0F78:q <= 8'h06;
            12'h0F79:q <= 8'h09;
            12'h0F7A:q <= 8'h10;
            12'h0F7B:q <= 8'h1E;
            12'h0F7C:q <= 8'h17;
            12'h0F7D:q <= 8'h1B;
            12'h0F7E:q <= 8'h24;
            12'h0F7F:q <= 8'h1E;
            12'h0F80:q <= 8'h12;
            12'h0F81:q <= 8'h12;
            12'h0F82:q <= 8'h00;
            12'h0F83:q <= 8'h10;
            12'h0F84:q <= 8'hFF;
            12'h0F85:q <= 8'h07;
            12'h0F86:q <= 8'h1F;
            12'h0F87:q <= 8'h03;
            12'h0F88:q <= 8'h12;
            12'h0F89:q <= 8'h27;
            12'h0F8A:q <= 8'h26;
            12'h0F8B:q <= 8'h22;
            12'h0F8C:q <= 8'h0F;
            12'h0F8D:q <= 8'h1A;
            12'h0F8E:q <= 8'h2C;
            12'h0F8F:q <= 8'h02;
            12'h0F90:q <= 8'h01;
            12'h0F91:q <= 8'hFF;
            12'h0F92:q <= 8'h08;
            12'h0F93:q <= 8'h16;
            12'h0F94:q <= 8'h29;
            12'h0F95:q <= 8'h0B;
            12'h0F96:q <= 8'h20;
            12'h0F97:q <= 8'h03;
            12'h0F98:q <= 8'h1B;
            12'h0F99:q <= 8'h14;
            12'h0F9A:q <= 8'h06;
            12'h0F9B:q <= 8'h19;
            12'h0F9C:q <= 8'h03;
            12'h0F9D:q <= 8'h08;
            12'h0F9E:q <= 8'hFF;
            12'h0F9F:q <= 8'h09;
            12'h0FA0:q <= 8'h25;
            12'h0FA1:q <= 8'h0A;
            12'h0FA2:q <= 8'h19;
            12'h0FA3:q <= 8'h06;
            12'h0FA4:q <= 8'h10;
            12'h0FA5:q <= 8'h01;
            12'h0FA6:q <= 8'h16;
            12'h0FA7:q <= 8'h18;
            12'h0FA8:q <= 8'h05;
            12'h0FA9:q <= 8'h1B;
            12'h0FAA:q <= 8'h07;
            12'h0FAB:q <= 8'hFF;
            12'h0FAC:q <= 8'h0A;
            12'h0FAD:q <= 8'h00;
            12'h0FAE:q <= 8'h08;
            12'h0FAF:q <= 8'h14;
            12'h0FB0:q <= 8'h04;
            12'h0FB1:q <= 8'h0F;
            12'h0FB2:q <= 8'h27;
            12'h0FB3:q <= 8'h21;
            12'h0FB4:q <= 8'h1C;
            12'h0FB5:q <= 8'h26;
            12'h0FB6:q <= 8'h1E;
            12'h0FB7:q <= 8'h0D;
            12'h0FB8:q <= 8'hFF;
            12'h0FB9:q <= 8'h0B;
            12'h0FBA:q <= 8'h0D;
            12'h0FBB:q <= 8'h12;
            12'h0FBC:q <= 8'h1D;
            12'h0FBD:q <= 8'h23;
            12'h0FBE:q <= 8'h2B;
            12'h0FBF:q <= 8'h15;
            12'h0FC0:q <= 8'h28;
            12'h0FC1:q <= 8'h19;
            12'h0FC2:q <= 8'h18;
            12'h0FC3:q <= 8'h29;
            12'h0FC4:q <= 8'h04;
            12'h0FC5:q <= 8'hFF;
            12'h0FC6:q <= 8'h0C;
            12'h0FC7:q <= 8'h0A;
            12'h0FC8:q <= 8'h06;
            12'h0FC9:q <= 8'h0C;
            12'h0FCA:q <= 8'h22;
            12'h0FCB:q <= 8'h2C;
            12'h0FCC:q <= 8'h13;
            12'h0FCD:q <= 8'h0E;
            12'h0FCE:q <= 8'h08;
            12'h0FCF:q <= 8'h28;
            12'h0FD0:q <= 8'h25;
            12'h0FD1:q <= 8'h1D;
            12'h0FD2:q <= 8'hFF;
            12'h0FD3:q <= 8'h0D;
            12'h0FD4:q <= 8'h24;
            12'h0FD5:q <= 8'h28;
            12'h0FD6:q <= 8'h0A;
            12'h0FD7:q <= 8'h0D;
            12'h0FD8:q <= 8'h07;
            12'h0FD9:q <= 8'h29;
            12'h0FDA:q <= 8'h25;
            12'h0FDB:q <= 8'h1F;
            12'h0FDC:q <= 8'h13;
            12'h0FDD:q <= 8'h0E;
            12'h0FDE:q <= 8'h0C;
            12'h0FDF:q <= 8'hFF;
            12'h0FE0:q <= 8'h0E;
            12'h0FE1:q <= 8'h12;
            12'h0FE2:q <= 8'h25;
            12'h0FE3:q <= 8'h1C;
            12'h0FE4:q <= 8'h1A;
            12'h0FE5:q <= 8'h21;
            12'h0FE6:q <= 8'h23;
            12'h0FE7:q <= 8'h26;
            12'h0FE8:q <= 8'h07;
            12'h0FE9:q <= 8'h1A;
            12'h0FEA:q <= 8'h21;
            12'h0FEB:q <= 8'h1C;
            12'h0FEC:q <= 8'hFF;
            12'h0FED:q <= 8'h0F;
            12'h0FEE:q <= 8'h2C;
            12'h0FEF:q <= 8'h0B;
            12'h0FF0:q <= 8'hFF;
            12'h0FF1:q <= 8'h10;
            12'h0FF2:q <= 8'h06;
            12'h0FF3:q <= 8'h15;
            12'h0FF4:q <= 8'hFF;
            12'h0FF5:q <= 8'h11;
            12'h0FF6:q <= 8'h03;
            12'h0FF7:q <= 8'h20;
            12'h0FF8:q <= 8'hFF;
            12'h0FF9:q <= 8'h12;
            12'h0FFA:q <= 8'h1D;
            12'h0FFB:q <= 8'h0F;
            12'h0FFC:q <= 8'hFF;
            12'h0FFD:q <= 8'h13;
            12'h0FFE:q <= 8'h07;
            12'h0FFF:q <= 8'h27;
            12'h1000:q <= 8'hFF;
            12'h1001:q <= 8'h14;
            12'h1002:q <= 8'h1B;
            12'h1003:q <= 8'h1E;
            12'h1004:q <= 8'hFF;
            12'h1005:q <= 8'h15;
            12'h1006:q <= 8'h08;
            12'h1007:q <= 8'h26;
            12'h1008:q <= 8'hFF;
            12'h1009:q <= 8'h16;
            12'h100A:q <= 8'h0E;
            12'h100B:q <= 8'h19;
            12'h100C:q <= 8'hFF;
            12'h100D:q <= 8'h17;
            12'h100E:q <= 8'h0B;
            12'h100F:q <= 8'h17;
            12'h1010:q <= 8'hFF;
            12'h1011:q <= 8'h18;
            12'h1012:q <= 8'h2A;
            12'h1013:q <= 8'h2A;
            12'h1014:q <= 8'hFF;
            12'h1015:q <= 8'h19;
            12'h1016:q <= 8'h1A;
            12'h1017:q <= 8'h1C;
            12'h1018:q <= 8'hFF;
            12'h1019:q <= 8'h1A;
            12'h101A:q <= 8'h0F;
            12'h101B:q <= 8'h23;
            12'h101C:q <= 8'hFF;
            12'h101D:q <= 8'h1B;
            12'h101E:q <= 8'h14;
            12'h101F:q <= 8'h18;
            12'h1020:q <= 8'hFF;
            12'h1021:q <= 8'h1C;
            12'h1022:q <= 8'h11;
            12'h1023:q <= 8'h24;
            12'h1024:q <= 8'hFF;
            12'h1025:q <= 8'h1D;
            12'h1026:q <= 8'h04;
            12'h1027:q <= 8'h09;
            12'h1028:q <= 8'hFF;
            12'h1029:q <= 8'h1E;
            12'h102A:q <= 8'h05;
            12'h102B:q <= 8'h02;
            12'h102C:q <= 8'hFF;
            12'h102D:q <= 8'h1F;
            12'h102E:q <= 8'h0C;
            12'h102F:q <= 8'h00;
            12'h1030:q <= 8'hFF;
            12'h1031:q <= 8'h20;
            12'h1032:q <= 8'h27;
            12'h1033:q <= 8'h05;
            12'h1034:q <= 8'hFF;
            12'h1035:q <= 8'h21;
            12'h1036:q <= 8'h26;
            12'h1037:q <= 8'h07;
            12'h1038:q <= 8'hFF;
            12'h1039:q <= 8'h22;
            12'h103A:q <= 8'h22;
            12'h103B:q <= 8'h1B;
            12'h103C:q <= 8'hFF;
            12'h103D:q <= 8'h23;
            12'h103E:q <= 8'h10;
            12'h103F:q <= 8'h13;
            12'h1040:q <= 8'hFF;
            12'h1041:q <= 8'h24;
            12'h1042:q <= 8'h17;
            12'h1043:q <= 8'h04;
            12'h1044:q <= 8'hFF;
            12'h1045:q <= 8'h25;
            12'h1046:q <= 8'h21;
            12'h1047:q <= 8'h22;
            12'h1048:q <= 8'hFF;
            12'h1049:q <= 8'h26;
            12'h104A:q <= 8'h18;
            12'h104B:q <= 8'h14;
            12'h104C:q <= 8'hFF;
            12'h104D:q <= 8'h27;
            12'h104E:q <= 8'h01;
            12'h104F:q <= 8'h11;
            12'h1050:q <= 8'hFF;
            12'h1051:q <= 8'h28;
            12'h1052:q <= 8'h02;
            12'h1053:q <= 8'h01;
            12'h1054:q <= 8'hFF;
            12'h1055:q <= 8'h29;
            12'h1056:q <= 8'h2B;
            12'h1057:q <= 8'h0D;
            12'h1058:q <= 8'hFF;
            12'h1059:q <= 8'h2A;
            12'h105A:q <= 8'h19;
            12'h105B:q <= 8'h21;
            12'h105C:q <= 8'hFF;
            12'h105D:q <= 8'h2B;
            12'h105E:q <= 8'h1C;
            12'h105F:q <= 8'h2C;
            12'h1060:q <= 8'hFF;
            12'h1061:q <= 8'h2C;
            12'h1062:q <= 8'h29;
            12'h1063:q <= 8'h1F;
            12'h1064:q <= 8'hFF;
            12'h1065:q <= 8'h00;
            12'h1066:q <= 8'h20;
            12'h1067:q <= 8'h04;
            12'h1068:q <= 8'hFF;
            12'h1069:q <= 8'h01;
            12'h106A:q <= 8'h04;
            12'h106B:q <= 8'h14;
            12'h106C:q <= 8'hFF;
            12'h106D:q <= 8'h02;
            12'h106E:q <= 8'h1B;
            12'h106F:q <= 8'h07;
            12'h1070:q <= 8'hFF;
            12'h1071:q <= 8'h03;
            12'h1072:q <= 8'h06;
            12'h1073:q <= 8'h03;
            12'h1074:q <= 8'hFF;
            12'h1075:q <= 8'h04;
            12'h1076:q <= 8'h27;
            12'h1077:q <= 8'h1D;
            12'h1078:q <= 8'hFF;
            12'h1079:q <= 8'h05;
            12'h107A:q <= 8'h03;
            12'h107B:q <= 8'h12;
            12'h107C:q <= 8'hFF;
            12'h107D:q <= 8'h06;
            12'h107E:q <= 8'h02;
            12'h107F:q <= 8'h0E;
            12'h1080:q <= 8'hFF;
            12'h1081:q <= 8'h07;
            12'h1082:q <= 8'h0C;
            12'h1083:q <= 8'h21;
            12'h1084:q <= 8'hFF;
            12'h1085:q <= 8'h08;
            12'h1086:q <= 8'h0D;
            12'h1087:q <= 8'h23;
            12'h1088:q <= 8'hFF;
            12'h1089:q <= 8'h09;
            12'h108A:q <= 8'h2A;
            12'h108B:q <= 8'h25;
            12'h108C:q <= 8'hFF;
            12'h108D:q <= 8'h0A;
            12'h108E:q <= 8'h17;
            12'h108F:q <= 8'h08;
            12'h1090:q <= 8'hFF;
            12'h1091:q <= 8'h0B;
            12'h1092:q <= 8'h15;
            12'h1093:q <= 8'h0B;
            12'h1094:q <= 8'hFF;
            12'h1095:q <= 8'h0C;
            12'h1096:q <= 8'h0B;
            12'h1097:q <= 8'h09;
            12'h1098:q <= 8'hFF;
            12'h1099:q <= 8'h0D;
            12'h109A:q <= 8'h22;
            12'h109B:q <= 8'h1A;
            12'h109C:q <= 8'hFF;
            12'h109D:q <= 8'h0E;
            12'h109E:q <= 8'h1F;
            12'h109F:q <= 8'h00;
            12'h10A0:q <= 8'hFF;
            12'h10A1:q <= 8'h0F;
            12'h10A2:q <= 8'h12;
            12'h10A3:q <= 8'h2C;
            12'h10A4:q <= 8'hFF;
            12'h10A5:q <= 8'h10;
            12'h10A6:q <= 8'h28;
            12'h10A7:q <= 8'h22;
            12'h10A8:q <= 8'hFF;
            12'h10A9:q <= 8'h11;
            12'h10AA:q <= 8'h0E;
            12'h10AB:q <= 8'h01;
            12'h10AC:q <= 8'hFF;
            12'h10AD:q <= 8'h12;
            12'h10AE:q <= 8'h0A;
            12'h10AF:q <= 8'h2A;
            12'h10B0:q <= 8'hFF;
            12'h10B1:q <= 8'h13;
            12'h10B2:q <= 8'h26;
            12'h10B3:q <= 8'h17;
            12'h10B4:q <= 8'hFF;
            12'h10B5:q <= 8'h14;
            12'h10B6:q <= 8'h21;
            12'h10B7:q <= 8'h1E;
            12'h10B8:q <= 8'hFF;
            12'h10B9:q <= 8'h15;
            12'h10BA:q <= 8'h07;
            12'h10BB:q <= 8'h24;
            12'h10BC:q <= 8'hFF;
            12'h10BD:q <= 8'h16;
            12'h10BE:q <= 8'h1A;
            12'h10BF:q <= 8'h28;
            12'h10C0:q <= 8'hFF;
            12'h10C1:q <= 8'h17;
            12'h10C2:q <= 8'h0F;
            12'h10C3:q <= 8'h0D;
            12'h10C4:q <= 8'hFF;
            12'h10C5:q <= 8'h18;
            12'h10C6:q <= 8'h00;
            12'h10C7:q <= 8'h11;
            12'h10C8:q <= 8'hFF;
            12'h10C9:q <= 8'h19;
            12'h10CA:q <= 8'h1E;
            12'h10CB:q <= 8'h20;
            12'h10CC:q <= 8'hFF;
            12'h10CD:q <= 8'h1A;
            12'h10CE:q <= 8'h1C;
            12'h10CF:q <= 8'h1F;
            12'h10D0:q <= 8'hFF;
            12'h10D1:q <= 8'h1B;
            12'h10D2:q <= 8'h2B;
            12'h10D3:q <= 8'h29;
            12'h10D4:q <= 8'hFF;
            12'h10D5:q <= 8'h1C;
            12'h10D6:q <= 8'h05;
            12'h10D7:q <= 8'h1B;
            12'h10D8:q <= 8'hFF;
            12'h10D9:q <= 8'h1D;
            12'h10DA:q <= 8'h14;
            12'h10DB:q <= 8'h2B;
            12'h10DC:q <= 8'hFF;
            12'h10DD:q <= 8'h1E;
            12'h10DE:q <= 8'h2C;
            12'h10DF:q <= 8'h1C;
            12'h10E0:q <= 8'hFF;
            12'h10E1:q <= 8'h1F;
            12'h10E2:q <= 8'h25;
            12'h10E3:q <= 8'h0C;
            12'h10E4:q <= 8'hFF;
            12'h10E5:q <= 8'h20;
            12'h10E6:q <= 8'h13;
            12'h10E7:q <= 8'h05;
            12'h10E8:q <= 8'hFF;
            12'h10E9:q <= 8'h21;
            12'h10EA:q <= 8'h18;
            12'h10EB:q <= 8'h0A;
            12'h10EC:q <= 8'hFF;
            12'h10ED:q <= 8'h22;
            12'h10EE:q <= 8'h24;
            12'h10EF:q <= 8'h19;
            12'h10F0:q <= 8'hFF;
            12'h10F1:q <= 8'h23;
            12'h10F2:q <= 8'h1D;
            12'h10F3:q <= 8'h18;
            12'h10F4:q <= 8'hFF;
            12'h10F5:q <= 8'h24;
            12'h10F6:q <= 8'h19;
            12'h10F7:q <= 8'h16;
            12'h10F8:q <= 8'hFF;
            12'h10F9:q <= 8'h25;
            12'h10FA:q <= 8'h01;
            12'h10FB:q <= 8'h15;
            12'h10FC:q <= 8'hFF;
            12'h10FD:q <= 8'h26;
            12'h10FE:q <= 8'h29;
            12'h10FF:q <= 8'h27;
            12'h1100:q <= 8'hFF;
            12'h1101:q <= 8'h27;
            12'h1102:q <= 8'h16;
            12'h1103:q <= 8'h10;
            12'h1104:q <= 8'hFF;
            12'h1105:q <= 8'h28;
            12'h1106:q <= 8'h10;
            12'h1107:q <= 8'h02;
            12'h1108:q <= 8'hFF;
            12'h1109:q <= 8'h29;
            12'h110A:q <= 8'h23;
            12'h110B:q <= 8'h0F;
            12'h110C:q <= 8'hFF;
            12'h110D:q <= 8'h2A;
            12'h110E:q <= 8'h09;
            12'h110F:q <= 8'h13;
            12'h1110:q <= 8'hFF;
            12'h1111:q <= 8'h2B;
            12'h1112:q <= 8'h11;
            12'h1113:q <= 8'h26;
            12'h1114:q <= 8'hFF;
            12'h1115:q <= 8'h2C;
            12'h1116:q <= 8'h08;
            12'h1117:q <= 8'h06;
            12'h1118:q <= 8'hFF;
            12'h1119:q <= 8'h00;
            12'h111A:q <= 8'h0C;
            12'h111B:q <= 8'h02;
            12'h111C:q <= 8'hFF;
            12'h111D:q <= 8'h01;
            12'h111E:q <= 8'h10;
            12'h111F:q <= 8'h1E;
            12'h1120:q <= 8'hFF;
            12'h1121:q <= 8'h02;
            12'h1122:q <= 8'h19;
            12'h1123:q <= 8'h1D;
            12'h1124:q <= 8'hFF;
            12'h1125:q <= 8'h03;
            12'h1126:q <= 8'h2C;
            12'h1127:q <= 8'h2A;
            12'h1128:q <= 8'hFF;
            12'h1129:q <= 8'h04;
            12'h112A:q <= 8'h00;
            12'h112B:q <= 8'h05;
            12'h112C:q <= 8'hFF;
            12'h112D:q <= 8'h05;
            12'h112E:q <= 8'h21;
            12'h112F:q <= 8'h29;
            12'h1130:q <= 8'hFF;
            12'h1131:q <= 8'h06;
            12'h1132:q <= 8'h13;
            12'h1133:q <= 8'h08;
            12'h1134:q <= 8'hFF;
            12'h1135:q <= 8'h07;
            12'h1136:q <= 8'h0B;
            12'h1137:q <= 8'h1B;
            12'h1138:q <= 8'hFF;
            12'h1139:q <= 8'h08;
            12'h113A:q <= 8'h06;
            12'h113B:q <= 8'h16;
            12'h113C:q <= 8'hFF;
            12'h113D:q <= 8'h09;
            12'h113E:q <= 8'h1F;
            12'h113F:q <= 8'h0A;
            12'h1140:q <= 8'hFF;
            12'h1141:q <= 8'h0A;
            12'h1142:q <= 8'h0A;
            12'h1143:q <= 8'h04;
            12'h1144:q <= 8'hFF;
            12'h1145:q <= 8'h0B;
            12'h1146:q <= 8'h25;
            12'h1147:q <= 8'h27;
            12'h1148:q <= 8'hFF;
            12'h1149:q <= 8'h0C;
            12'h114A:q <= 8'h11;
            12'h114B:q <= 8'h0F;
            12'h114C:q <= 8'hFF;
            12'h114D:q <= 8'h0D;
            12'h114E:q <= 8'h15;
            12'h114F:q <= 8'h28;
            12'h1150:q <= 8'hFF;
            12'h1151:q <= 8'h0E;
            12'h1152:q <= 8'h1D;
            12'h1153:q <= 8'h0C;
            12'h1154:q <= 8'hFF;
            12'h1155:q <= 8'h0F;
            12'h1156:q <= 8'h0E;
            12'h1157:q <= 8'h22;
            12'h1158:q <= 8'hFF;
            12'h1159:q <= 8'h10;
            12'h115A:q <= 8'h17;
            12'h115B:q <= 8'h06;
            12'h115C:q <= 8'hFF;
            12'h115D:q <= 8'h11;
            12'h115E:q <= 8'h04;
            12'h115F:q <= 8'h0D;
            12'h1160:q <= 8'hFF;
            12'h1161:q <= 8'h12;
            12'h1162:q <= 8'h09;
            12'h1163:q <= 8'h07;
            12'h1164:q <= 8'hFF;
            12'h1165:q <= 8'h13;
            12'h1166:q <= 8'h22;
            12'h1167:q <= 8'h17;
            12'h1168:q <= 8'hFF;
            12'h1169:q <= 8'h14;
            12'h116A:q <= 8'h0D;
            12'h116B:q <= 8'h15;
            12'h116C:q <= 8'hFF;
            12'h116D:q <= 8'h15;
            12'h116E:q <= 8'h27;
            12'h116F:q <= 8'h09;
            12'h1170:q <= 8'hFF;
            12'h1171:q <= 8'h16;
            12'h1172:q <= 8'h1C;
            12'h1173:q <= 8'h23;
            12'h1174:q <= 8'hFF;
            12'h1175:q <= 8'h17;
            12'h1176:q <= 8'h14;
            12'h1177:q <= 8'h01;
            12'h1178:q <= 8'hFF;
            12'h1179:q <= 8'h18;
            12'h117A:q <= 8'h02;
            12'h117B:q <= 8'h10;
            12'h117C:q <= 8'hFF;
            12'h117D:q <= 8'h19;
            12'h117E:q <= 8'h2B;
            12'h117F:q <= 8'h2B;
            12'h1180:q <= 8'hFF;
            12'h1181:q <= 8'h1A;
            12'h1182:q <= 8'h08;
            12'h1183:q <= 8'h0E;
            12'h1184:q <= 8'hFF;
            12'h1185:q <= 8'h1B;
            12'h1186:q <= 8'h2A;
            12'h1187:q <= 8'h24;
            12'h1188:q <= 8'hFF;
            12'h1189:q <= 8'h1C;
            12'h118A:q <= 8'h1B;
            12'h118B:q <= 8'h19;
            12'h118C:q <= 8'hFF;
            12'h118D:q <= 8'h1D;
            12'h118E:q <= 8'h12;
            12'h118F:q <= 8'h20;
            12'h1190:q <= 8'hFF;
            12'h1191:q <= 8'h1E;
            12'h1192:q <= 8'h16;
            12'h1193:q <= 8'h1A;
            12'h1194:q <= 8'hFF;
            12'h1195:q <= 8'h1F;
            12'h1196:q <= 8'h28;
            12'h1197:q <= 8'h12;
            12'h1198:q <= 8'hFF;
            12'h1199:q <= 8'h20;
            12'h119A:q <= 8'h23;
            12'h119B:q <= 8'h0B;
            12'h119C:q <= 8'hFF;
            12'h119D:q <= 8'h21;
            12'h119E:q <= 8'h07;
            12'h119F:q <= 8'h03;
            12'h11A0:q <= 8'hFF;
            12'h11A1:q <= 8'h22;
            12'h11A2:q <= 8'h24;
            12'h11A3:q <= 8'h18;
            12'h11A4:q <= 8'hFF;
            12'h11A5:q <= 8'h23;
            12'h11A6:q <= 8'h0F;
            12'h11A7:q <= 8'h26;
            12'h11A8:q <= 8'hFF;
            12'h11A9:q <= 8'h24;
            12'h11AA:q <= 8'h1E;
            12'h11AB:q <= 8'h00;
            12'h11AC:q <= 8'hFF;
            12'h11AD:q <= 8'h25;
            12'h11AE:q <= 8'h20;
            12'h11AF:q <= 8'h13;
            12'h11B0:q <= 8'hFF;
            12'h11B1:q <= 8'h26;
            12'h11B2:q <= 8'h1A;
            12'h11B3:q <= 8'h1C;
            12'h11B4:q <= 8'hFF;
            12'h11B5:q <= 8'h27;
            12'h11B6:q <= 8'h01;
            12'h11B7:q <= 8'h11;
            12'h11B8:q <= 8'hFF;
            12'h11B9:q <= 8'h28;
            12'h11BA:q <= 8'h26;
            12'h11BB:q <= 8'h21;
            12'h11BC:q <= 8'hFF;
            12'h11BD:q <= 8'h29;
            12'h11BE:q <= 8'h05;
            12'h11BF:q <= 8'h2C;
            12'h11C0:q <= 8'hFF;
            12'h11C1:q <= 8'h2A;
            12'h11C2:q <= 8'h29;
            12'h11C3:q <= 8'h14;
            12'h11C4:q <= 8'hFF;
            12'h11C5:q <= 8'h2B;
            12'h11C6:q <= 8'h18;
            12'h11C7:q <= 8'h25;
            12'h11C8:q <= 8'hFF;
            12'h11C9:q <= 8'h2C;
            12'h11CA:q <= 8'h03;
            12'h11CB:q <= 8'h1F;
            12'h11CC:q <= 8'hFF;
            12'h11CD:q <= 8'h03;
            12'h11CE:q <= 8'h06;
            12'h11CF:q <= 8'h0A;
            12'h11D0:q <= 8'h07;
            12'h11D1:q <= 8'h05;
            12'h11D2:q <= 8'h01;
            12'h11D3:q <= 8'h00;
            12'h11D4:q <= 8'h04;
            12'h11D5:q <= 8'h05;
            12'h11D6:q <= 8'h02;
            12'h11D7:q <= 8'h0B;
            12'h11D8:q <= 8'h01;
            12'h11D9:q <= 8'hFF;
            12'h11DA:q <= 8'h04;
            12'h11DB:q <= 8'h05;
            12'h11DC:q <= 8'h0B;
            12'h11DD:q <= 8'hFF;
            12'h11DE:q <= 8'h05;
            12'h11DF:q <= 8'h0B;
            12'h11E0:q <= 8'h07;
            12'h11E1:q <= 8'hFF;
            12'h11E2:q <= 8'h06;
            12'h11E3:q <= 8'h09;
            12'h11E4:q <= 8'h01;
            12'h11E5:q <= 8'hFF;
            12'h11E6:q <= 8'h07;
            12'h11E7:q <= 8'h02;
            12'h11E8:q <= 8'h05;
            12'h11E9:q <= 8'hFF;
            12'h11EA:q <= 8'h08;
            12'h11EB:q <= 8'h01;
            12'h11EC:q <= 8'h08;
            12'h11ED:q <= 8'hFF;
            12'h11EE:q <= 8'h09;
            12'h11EF:q <= 8'h08;
            12'h11F0:q <= 8'h06;
            12'h11F1:q <= 8'hFF;
            12'h11F2:q <= 8'h0A;
            12'h11F3:q <= 8'h0A;
            12'h11F4:q <= 8'h02;
            12'h11F5:q <= 8'hFF;
            12'h11F6:q <= 8'h0B;
            12'h11F7:q <= 8'h07;
            12'h11F8:q <= 8'h00;
            12'h11F9:q <= 8'hFF;
            12'h11FA:q <= 8'h00;
            12'h11FB:q <= 8'h06;
            12'h11FC:q <= 8'h07;
            12'h11FD:q <= 8'hFF;
            12'h11FE:q <= 8'h01;
            12'h11FF:q <= 8'h03;
            12'h1200:q <= 8'h08;
            12'h1201:q <= 8'hFF;
            12'h1202:q <= 8'h02;
            12'h1203:q <= 8'h09;
            12'h1204:q <= 8'h00;
            12'h1205:q <= 8'hFF;
            12'h1206:q <= 8'h03;
            12'h1207:q <= 8'h00;
            12'h1208:q <= 8'h05;
            12'h1209:q <= 8'hFF;
            12'h120A:q <= 8'h04;
            12'h120B:q <= 8'h05;
            12'h120C:q <= 8'h02;
            12'h120D:q <= 8'hFF;
            12'h120E:q <= 8'h05;
            12'h120F:q <= 8'h0A;
            12'h1210:q <= 8'h03;
            12'h1211:q <= 8'hFF;
            12'h1212:q <= 8'h06;
            12'h1213:q <= 8'h08;
            12'h1214:q <= 8'h09;
            12'h1215:q <= 8'hFF;
            12'h1216:q <= 8'h07;
            12'h1217:q <= 8'h02;
            12'h1218:q <= 8'h0A;
            12'h1219:q <= 8'hFF;
            12'h121A:q <= 8'h08;
            12'h121B:q <= 8'h07;
            12'h121C:q <= 8'h01;
            12'h121D:q <= 8'hFF;
            12'h121E:q <= 8'h09;
            12'h121F:q <= 8'h04;
            12'h1220:q <= 8'h04;
            12'h1221:q <= 8'hFF;
            12'h1222:q <= 8'h0A;
            12'h1223:q <= 8'h0B;
            12'h1224:q <= 8'h06;
            12'h1225:q <= 8'hFF;
            12'h1226:q <= 8'h0B;
            12'h1227:q <= 8'h01;
            12'h1228:q <= 8'h0B;
            12'h1229:q <= 8'hFF;
            12'h122A:q <= 8'h00;
            12'h122B:q <= 8'h08;
            12'h122C:q <= 8'h07;
            12'h122D:q <= 8'hFF;
            12'h122E:q <= 8'h01;
            12'h122F:q <= 8'h09;
            12'h1230:q <= 8'h08;
            12'h1231:q <= 8'hFF;
            12'h1232:q <= 8'h02;
            12'h1233:q <= 8'h05;
            12'h1234:q <= 8'h0B;
            12'h1235:q <= 8'hFF;
            12'h1236:q <= 8'h03;
            12'h1237:q <= 8'h01;
            12'h1238:q <= 8'h03;
            12'h1239:q <= 8'hFF;
            12'h123A:q <= 8'h04;
            12'h123B:q <= 8'h07;
            12'h123C:q <= 8'h01;
            12'h123D:q <= 8'hFF;
            12'h123E:q <= 8'h05;
            12'h123F:q <= 8'h06;
            12'h1240:q <= 8'h02;
            12'h1241:q <= 8'hFF;
            12'h1242:q <= 8'h06;
            12'h1243:q <= 8'h00;
            12'h1244:q <= 8'h0A;
            12'h1245:q <= 8'hFF;
            12'h1246:q <= 8'h07;
            12'h1247:q <= 8'h0A;
            12'h1248:q <= 8'h05;
            12'h1249:q <= 8'hFF;
            12'h124A:q <= 8'h08;
            12'h124B:q <= 8'h02;
            12'h124C:q <= 8'h09;
            12'h124D:q <= 8'hFF;
            12'h124E:q <= 8'h09;
            12'h124F:q <= 8'h03;
            12'h1250:q <= 8'h06;
            12'h1251:q <= 8'hFF;
            12'h1252:q <= 8'h0A;
            12'h1253:q <= 8'h04;
            12'h1254:q <= 8'h04;
            12'h1255:q <= 8'hFF;
            12'h1256:q <= 8'h0B;
            12'h1257:q <= 8'h0B;
            12'h1258:q <= 8'h00;
            12'h1259:q <= 8'hFF;
            12'h125A:q <= 8'h00;
            12'h125B:q <= 8'h05;
            12'h125C:q <= 8'h10;
            12'h125D:q <= 8'h1F;
            12'h125E:q <= 8'h18;
            12'h125F:q <= 8'h1F;
            12'h1260:q <= 8'h08;
            12'h1261:q <= 8'h09;
            12'h1262:q <= 8'h0C;
            12'h1263:q <= 8'h12;
            12'h1264:q <= 8'h0C;
            12'h1265:q <= 8'hFF;
            12'h1266:q <= 8'h01;
            12'h1267:q <= 8'h11;
            12'h1268:q <= 8'h16;
            12'h1269:q <= 8'h15;
            12'h126A:q <= 8'h1E;
            12'h126B:q <= 8'h11;
            12'h126C:q <= 8'h1A;
            12'h126D:q <= 8'h20;
            12'h126E:q <= 8'h11;
            12'h126F:q <= 8'h23;
            12'h1270:q <= 8'h09;
            12'h1271:q <= 8'hFF;
            12'h1272:q <= 8'h02;
            12'h1273:q <= 8'h1E;
            12'h1274:q <= 8'h09;
            12'h1275:q <= 8'h0C;
            12'h1276:q <= 8'h1D;
            12'h1277:q <= 8'h14;
            12'h1278:q <= 8'h09;
            12'h1279:q <= 8'h18;
            12'h127A:q <= 8'h13;
            12'h127B:q <= 8'h14;
            12'h127C:q <= 8'h21;
            12'h127D:q <= 8'hFF;
            12'h127E:q <= 8'h03;
            12'h127F:q <= 8'h23;
            12'h1280:q <= 8'h14;
            12'h1281:q <= 8'h22;
            12'h1282:q <= 8'h1C;
            12'h1283:q <= 8'h21;
            12'h1284:q <= 8'h0A;
            12'h1285:q <= 8'h0F;
            12'h1286:q <= 8'h19;
            12'h1287:q <= 8'h0D;
            12'h1288:q <= 8'h1C;
            12'h1289:q <= 8'hFF;
            12'h128A:q <= 8'h04;
            12'h128B:q <= 8'h07;
            12'h128C:q <= 8'h13;
            12'h128D:q <= 8'h04;
            12'h128E:q <= 8'h17;
            12'h128F:q <= 8'h23;
            12'h1290:q <= 8'h0D;
            12'h1291:q <= 8'h21;
            12'h1292:q <= 8'h0A;
            12'h1293:q <= 8'h22;
            12'h1294:q <= 8'h17;
            12'h1295:q <= 8'hFF;
            12'h1296:q <= 8'h05;
            12'h1297:q <= 8'h18;
            12'h1298:q <= 8'h0F;
            12'h1299:q <= 8'h03;
            12'h129A:q <= 8'h10;
            12'h129B:q <= 8'h13;
            12'h129C:q <= 8'h18;
            12'h129D:q <= 8'h1C;
            12'h129E:q <= 8'h05;
            12'h129F:q <= 8'h03;
            12'h12A0:q <= 8'h02;
            12'h12A1:q <= 8'hFF;
            12'h12A2:q <= 8'h06;
            12'h12A3:q <= 8'h1B;
            12'h12A4:q <= 8'h1C;
            12'h12A5:q <= 8'h16;
            12'h12A6:q <= 8'h1A;
            12'h12A7:q <= 8'h10;
            12'h12A8:q <= 8'h04;
            12'h12A9:q <= 8'h00;
            12'h12AA:q <= 8'h07;
            12'h12AB:q <= 8'h16;
            12'h12AC:q <= 8'h11;
            12'h12AD:q <= 8'hFF;
            12'h12AE:q <= 8'h07;
            12'h12AF:q <= 8'h0D;
            12'h12B0:q <= 8'h17;
            12'h12B1:q <= 8'h02;
            12'h12B2:q <= 8'h0E;
            12'h12B3:q <= 8'h0F;
            12'h12B4:q <= 8'h17;
            12'h12B5:q <= 8'h06;
            12'h12B6:q <= 8'h17;
            12'h12B7:q <= 8'h0F;
            12'h12B8:q <= 8'h04;
            12'h12B9:q <= 8'hFF;
            12'h12BA:q <= 8'h08;
            12'h12BB:q <= 8'h06;
            12'h12BC:q <= 8'h0B;
            12'h12BD:q <= 8'h08;
            12'h12BE:q <= 8'h11;
            12'h12BF:q <= 8'h1B;
            12'h12C0:q <= 8'h1E;
            12'h12C1:q <= 8'h1F;
            12'h12C2:q <= 8'h12;
            12'h12C3:q <= 8'h0B;
            12'h12C4:q <= 8'h20;
            12'h12C5:q <= 8'hFF;
            12'h12C6:q <= 8'h09;
            12'h12C7:q <= 8'h21;
            12'h12C8:q <= 8'h12;
            12'h12C9:q <= 8'h0D;
            12'h12CA:q <= 8'h05;
            12'h12CB:q <= 8'h03;
            12'h12CC:q <= 8'h01;
            12'h12CD:q <= 8'h1B;
            12'h12CE:q <= 8'h22;
            12'h12CF:q <= 8'h1A;
            12'h12D0:q <= 8'h08;
            12'h12D1:q <= 8'hFF;
            12'h12D2:q <= 8'h0A;
            12'h12D3:q <= 8'h0C;
            12'h12D4:q <= 8'h08;
            12'h12D5:q <= 8'h07;
            12'h12D6:q <= 8'h23;
            12'h12D7:q <= 8'h07;
            12'h12D8:q <= 8'h22;
            12'h12D9:q <= 8'h1A;
            12'h12DA:q <= 8'h02;
            12'h12DB:q <= 8'h1B;
            12'h12DC:q <= 8'h01;
            12'h12DD:q <= 8'hFF;
            12'h12DE:q <= 8'h0B;
            12'h12DF:q <= 8'h10;
            12'h12E0:q <= 8'h18;
            12'h12E1:q <= 8'h0F;
            12'h12E2:q <= 8'h20;
            12'h12E3:q <= 8'h06;
            12'h12E4:q <= 8'h0C;
            12'h12E5:q <= 8'h03;
            12'h12E6:q <= 8'h0E;
            12'h12E7:q <= 8'h06;
            12'h12E8:q <= 8'h13;
            12'h12E9:q <= 8'hFF;
            12'h12EA:q <= 8'h0C;
            12'h12EB:q <= 8'h0F;
            12'h12EC:q <= 8'h0A;
            12'h12ED:q <= 8'h21;
            12'h12EE:q <= 8'h0A;
            12'h12EF:q <= 8'h12;
            12'h12F0:q <= 8'h02;
            12'h12F1:q <= 8'h23;
            12'h12F2:q <= 8'h0B;
            12'h12F3:q <= 8'h1D;
            12'h12F4:q <= 8'h00;
            12'h12F5:q <= 8'hFF;
            12'h12F6:q <= 8'h0D;
            12'h12F7:q <= 8'h1A;
            12'h12F8:q <= 8'h1B;
            12'h12F9:q <= 8'h06;
            12'h12FA:q <= 8'h09;
            12'h12FB:q <= 8'h19;
            12'h12FC:q <= 8'h05;
            12'h12FD:q <= 8'h1D;
            12'h12FE:q <= 8'h15;
            12'h12FF:q <= 8'h0A;
            12'h1300:q <= 8'h1F;
            12'h1301:q <= 8'hFF;
            12'h1302:q <= 8'h0E;
            12'h1303:q <= 8'h1D;
            12'h1304:q <= 8'h19;
            12'h1305:q <= 8'h14;
            12'h1306:q <= 8'h01;
            12'h1307:q <= 8'h20;
            12'h1308:q <= 8'h15;
            12'h1309:q <= 8'h08;
            12'h130A:q <= 8'h1E;
            12'h130B:q <= 8'h07;
            12'h130C:q <= 8'h15;
            12'h130D:q <= 8'hFF;
            12'h130E:q <= 8'h0F;
            12'h130F:q <= 8'h00;
            12'h1310:q <= 8'h03;
            12'h1311:q <= 8'h1B;
            12'h1312:q <= 8'h0B;
            12'h1313:q <= 8'h00;
            12'h1314:q <= 8'h0B;
            12'h1315:q <= 8'h10;
            12'h1316:q <= 8'h04;
            12'h1317:q <= 8'h0E;
            12'h1318:q <= 8'h18;
            12'h1319:q <= 8'hFF;
            12'h131A:q <= 8'h10;
            12'h131B:q <= 8'h16;
            12'h131C:q <= 8'h21;
            12'h131D:q <= 8'h13;
            12'h131E:q <= 8'h12;
            12'h131F:q <= 8'h1D;
            12'h1320:q <= 8'h16;
            12'h1321:q <= 8'h16;
            12'h1322:q <= 8'h0D;
            12'h1323:q <= 8'h1E;
            12'h1324:q <= 8'h05;
            12'h1325:q <= 8'hFF;
            12'h1326:q <= 8'h11;
            12'h1327:q <= 8'h15;
            12'h1328:q <= 8'h11;
            12'h1329:q <= 8'h00;
            12'h132A:q <= 8'h19;
            12'h132B:q <= 8'h1C;
            12'h132C:q <= 8'h0E;
            12'h132D:q <= 8'h01;
            12'h132E:q <= 8'h14;
            12'h132F:q <= 8'h10;
            12'h1330:q <= 8'h19;
            12'h1331:q <= 8'hFF;
            12'h1332:q <= 8'h12;
            12'h1333:q <= 8'h03;
            12'h1334:q <= 8'h22;
            12'h1335:q <= 8'hFF;
            12'h1336:q <= 8'h13;
            12'h1337:q <= 8'h02;
            12'h1338:q <= 8'h07;
            12'h1339:q <= 8'hFF;
            12'h133A:q <= 8'h14;
            12'h133B:q <= 8'h08;
            12'h133C:q <= 8'h1A;
            12'h133D:q <= 8'hFF;
            12'h133E:q <= 8'h15;
            12'h133F:q <= 8'h13;
            12'h1340:q <= 8'h02;
            12'h1341:q <= 8'hFF;
            12'h1342:q <= 8'h16;
            12'h1343:q <= 8'h0E;
            12'h1344:q <= 8'h05;
            12'h1345:q <= 8'hFF;
            12'h1346:q <= 8'h17;
            12'h1347:q <= 8'h1F;
            12'h1348:q <= 8'h23;
            12'h1349:q <= 8'hFF;
            12'h134A:q <= 8'h18;
            12'h134B:q <= 8'h1C;
            12'h134C:q <= 8'h20;
            12'h134D:q <= 8'hFF;
            12'h134E:q <= 8'h19;
            12'h134F:q <= 8'h0A;
            12'h1350:q <= 8'h00;
            12'h1351:q <= 8'hFF;
            12'h1352:q <= 8'h1A;
            12'h1353:q <= 8'h09;
            12'h1354:q <= 8'h15;
            12'h1355:q <= 8'hFF;
            12'h1356:q <= 8'h1B;
            12'h1357:q <= 8'h01;
            12'h1358:q <= 8'h06;
            12'h1359:q <= 8'hFF;
            12'h135A:q <= 8'h1C;
            12'h135B:q <= 8'h19;
            12'h135C:q <= 8'h1D;
            12'h135D:q <= 8'hFF;
            12'h135E:q <= 8'h1D;
            12'h135F:q <= 8'h14;
            12'h1360:q <= 8'h0D;
            12'h1361:q <= 8'hFF;
            12'h1362:q <= 8'h1E;
            12'h1363:q <= 8'h04;
            12'h1364:q <= 8'h0C;
            12'h1365:q <= 8'hFF;
            12'h1366:q <= 8'h1F;
            12'h1367:q <= 8'h20;
            12'h1368:q <= 8'h04;
            12'h1369:q <= 8'hFF;
            12'h136A:q <= 8'h20;
            12'h136B:q <= 8'h22;
            12'h136C:q <= 8'h0E;
            12'h136D:q <= 8'hFF;
            12'h136E:q <= 8'h21;
            12'h136F:q <= 8'h0B;
            12'h1370:q <= 8'h01;
            12'h1371:q <= 8'hFF;
            12'h1372:q <= 8'h22;
            12'h1373:q <= 8'h17;
            12'h1374:q <= 8'h1F;
            12'h1375:q <= 8'hFF;
            12'h1376:q <= 8'h23;
            12'h1377:q <= 8'h12;
            12'h1378:q <= 8'h1E;
            12'h1379:q <= 8'hFF;
            12'h137A:q <= 8'h00;
            12'h137B:q <= 8'h09;
            12'h137C:q <= 8'h21;
            12'h137D:q <= 8'hFF;
            12'h137E:q <= 8'h01;
            12'h137F:q <= 8'h22;
            12'h1380:q <= 8'h1F;
            12'h1381:q <= 8'hFF;
            12'h1382:q <= 8'h02;
            12'h1383:q <= 8'h23;
            12'h1384:q <= 8'h13;
            12'h1385:q <= 8'hFF;
            12'h1386:q <= 8'h03;
            12'h1387:q <= 8'h00;
            12'h1388:q <= 8'h14;
            12'h1389:q <= 8'hFF;
            12'h138A:q <= 8'h04;
            12'h138B:q <= 8'h03;
            12'h138C:q <= 8'h1A;
            12'h138D:q <= 8'hFF;
            12'h138E:q <= 8'h05;
            12'h138F:q <= 8'h01;
            12'h1390:q <= 8'h1C;
            12'h1391:q <= 8'hFF;
            12'h1392:q <= 8'h06;
            12'h1393:q <= 8'h17;
            12'h1394:q <= 8'h06;
            12'h1395:q <= 8'hFF;
            12'h1396:q <= 8'h07;
            12'h1397:q <= 8'h20;
            12'h1398:q <= 8'h16;
            12'h1399:q <= 8'hFF;
            12'h139A:q <= 8'h08;
            12'h139B:q <= 8'h1B;
            12'h139C:q <= 8'h05;
            12'h139D:q <= 8'hFF;
            12'h139E:q <= 8'h09;
            12'h139F:q <= 8'h16;
            12'h13A0:q <= 8'h07;
            12'h13A1:q <= 8'hFF;
            12'h13A2:q <= 8'h0A;
            12'h13A3:q <= 8'h11;
            12'h13A4:q <= 8'h0C;
            12'h13A5:q <= 8'hFF;
            12'h13A6:q <= 8'h0B;
            12'h13A7:q <= 8'h1E;
            12'h13A8:q <= 8'h0A;
            12'h13A9:q <= 8'hFF;
            12'h13AA:q <= 8'h0C;
            12'h13AB:q <= 8'h02;
            12'h13AC:q <= 8'h20;
            12'h13AD:q <= 8'hFF;
            12'h13AE:q <= 8'h0D;
            12'h13AF:q <= 8'h04;
            12'h13B0:q <= 8'h00;
            12'h13B1:q <= 8'hFF;
            12'h13B2:q <= 8'h0E;
            12'h13B3:q <= 8'h1A;
            12'h13B4:q <= 8'h18;
            12'h13B5:q <= 8'hFF;
            12'h13B6:q <= 8'h0F;
            12'h13B7:q <= 8'h05;
            12'h13B8:q <= 8'h1E;
            12'h13B9:q <= 8'hFF;
            12'h13BA:q <= 8'h10;
            12'h13BB:q <= 8'h14;
            12'h13BC:q <= 8'h08;
            12'h13BD:q <= 8'hFF;
            12'h13BE:q <= 8'h11;
            12'h13BF:q <= 8'h1D;
            12'h13C0:q <= 8'h12;
            12'h13C1:q <= 8'hFF;
            12'h13C2:q <= 8'h12;
            12'h13C3:q <= 8'h13;
            12'h13C4:q <= 8'h04;
            12'h13C5:q <= 8'hFF;
            12'h13C6:q <= 8'h13;
            12'h13C7:q <= 8'h18;
            12'h13C8:q <= 8'h1D;
            12'h13C9:q <= 8'hFF;
            12'h13CA:q <= 8'h14;
            12'h13CB:q <= 8'h0B;
            12'h13CC:q <= 8'h15;
            12'h13CD:q <= 8'hFF;
            12'h13CE:q <= 8'h15;
            12'h13CF:q <= 8'h06;
            12'h13D0:q <= 8'h0F;
            12'h13D1:q <= 8'hFF;
            12'h13D2:q <= 8'h16;
            12'h13D3:q <= 8'h1C;
            12'h13D4:q <= 8'h03;
            12'h13D5:q <= 8'hFF;
            12'h13D6:q <= 8'h17;
            12'h13D7:q <= 8'h12;
            12'h13D8:q <= 8'h22;
            12'h13D9:q <= 8'hFF;
            12'h13DA:q <= 8'h18;
            12'h13DB:q <= 8'h15;
            12'h13DC:q <= 8'h09;
            12'h13DD:q <= 8'hFF;
            12'h13DE:q <= 8'h19;
            12'h13DF:q <= 8'h0C;
            12'h13E0:q <= 8'h17;
            12'h13E1:q <= 8'hFF;
            12'h13E2:q <= 8'h1A;
            12'h13E3:q <= 8'h10;
            12'h13E4:q <= 8'h0E;
            12'h13E5:q <= 8'hFF;
            12'h13E6:q <= 8'h1B;
            12'h13E7:q <= 8'h07;
            12'h13E8:q <= 8'h01;
            12'h13E9:q <= 8'hFF;
            12'h13EA:q <= 8'h1C;
            12'h13EB:q <= 8'h19;
            12'h13EC:q <= 8'h19;
            12'h13ED:q <= 8'hFF;
            12'h13EE:q <= 8'h1D;
            12'h13EF:q <= 8'h0A;
            12'h13F0:q <= 8'h0B;
            12'h13F1:q <= 8'hFF;
            12'h13F2:q <= 8'h1E;
            12'h13F3:q <= 8'h21;
            12'h13F4:q <= 8'h1B;
            12'h13F5:q <= 8'hFF;
            12'h13F6:q <= 8'h1F;
            12'h13F7:q <= 8'h0D;
            12'h13F8:q <= 8'h02;
            12'h13F9:q <= 8'hFF;
            12'h13FA:q <= 8'h20;
            12'h13FB:q <= 8'h0F;
            12'h13FC:q <= 8'h11;
            12'h13FD:q <= 8'hFF;
            12'h13FE:q <= 8'h21;
            12'h13FF:q <= 8'h0E;
            12'h1400:q <= 8'h10;
            12'h1401:q <= 8'hFF;
            12'h1402:q <= 8'h22;
            12'h1403:q <= 8'h08;
            12'h1404:q <= 8'h0D;
            12'h1405:q <= 8'hFF;
            12'h1406:q <= 8'h23;
            12'h1407:q <= 8'h1F;
            12'h1408:q <= 8'h23;
            12'h1409:q <= 8'hFF;
            12'h140A:q <= 8'h00;
            12'h140B:q <= 8'h1F;
            12'h140C:q <= 8'h03;
            12'h140D:q <= 8'hFF;
            12'h140E:q <= 8'h01;
            12'h140F:q <= 8'h07;
            12'h1410:q <= 8'h22;
            12'h1411:q <= 8'hFF;
            12'h1412:q <= 8'h02;
            12'h1413:q <= 8'h18;
            12'h1414:q <= 8'h1A;
            12'h1415:q <= 8'hFF;
            12'h1416:q <= 8'h03;
            12'h1417:q <= 8'h16;
            12'h1418:q <= 8'h0B;
            12'h1419:q <= 8'hFF;
            12'h141A:q <= 8'h04;
            12'h141B:q <= 8'h0D;
            12'h141C:q <= 8'h16;
            12'h141D:q <= 8'hFF;
            12'h141E:q <= 8'h05;
            12'h141F:q <= 8'h08;
            12'h1420:q <= 8'h15;
            12'h1421:q <= 8'hFF;
            12'h1422:q <= 8'h06;
            12'h1423:q <= 8'h02;
            12'h1424:q <= 8'h10;
            12'h1425:q <= 8'hFF;
            12'h1426:q <= 8'h07;
            12'h1427:q <= 8'h11;
            12'h1428:q <= 8'h14;
            12'h1429:q <= 8'hFF;
            12'h142A:q <= 8'h08;
            12'h142B:q <= 8'h0C;
            12'h142C:q <= 8'h1F;
            12'h142D:q <= 8'hFF;
            12'h142E:q <= 8'h09;
            12'h142F:q <= 8'h0A;
            12'h1430:q <= 8'h00;
            12'h1431:q <= 8'hFF;
            12'h1432:q <= 8'h0A;
            12'h1433:q <= 8'h13;
            12'h1434:q <= 8'h20;
            12'h1435:q <= 8'hFF;
            12'h1436:q <= 8'h0B;
            12'h1437:q <= 8'h0E;
            12'h1438:q <= 8'h0D;
            12'h1439:q <= 8'hFF;
            12'h143A:q <= 8'h0C;
            12'h143B:q <= 8'h22;
            12'h143C:q <= 8'h04;
            12'h143D:q <= 8'hFF;
            12'h143E:q <= 8'h0D;
            12'h143F:q <= 8'h1B;
            12'h1440:q <= 8'h0C;
            12'h1441:q <= 8'hFF;
            12'h1442:q <= 8'h0E;
            12'h1443:q <= 8'h00;
            12'h1444:q <= 8'h07;
            12'h1445:q <= 8'hFF;
            12'h1446:q <= 8'h0F;
            12'h1447:q <= 8'h1A;
            12'h1448:q <= 8'h0E;
            12'h1449:q <= 8'hFF;
            12'h144A:q <= 8'h10;
            12'h144B:q <= 8'h06;
            12'h144C:q <= 8'h06;
            12'h144D:q <= 8'hFF;
            12'h144E:q <= 8'h11;
            12'h144F:q <= 8'h17;
            12'h1450:q <= 8'h1D;
            12'h1451:q <= 8'hFF;
            12'h1452:q <= 8'h12;
            12'h1453:q <= 8'h0B;
            12'h1454:q <= 8'h1B;
            12'h1455:q <= 8'hFF;
            12'h1456:q <= 8'h13;
            12'h1457:q <= 8'h20;
            12'h1458:q <= 8'h23;
            12'h1459:q <= 8'hFF;
            12'h145A:q <= 8'h14;
            12'h145B:q <= 8'h15;
            12'h145C:q <= 8'h0A;
            12'h145D:q <= 8'hFF;
            12'h145E:q <= 8'h15;
            12'h145F:q <= 8'h12;
            12'h1460:q <= 8'h1C;
            12'h1461:q <= 8'hFF;
            12'h1462:q <= 8'h16;
            12'h1463:q <= 8'h03;
            12'h1464:q <= 8'h1E;
            12'h1465:q <= 8'hFF;
            12'h1466:q <= 8'h17;
            12'h1467:q <= 8'h19;
            12'h1468:q <= 8'h21;
            12'h1469:q <= 8'hFF;
            12'h146A:q <= 8'h18;
            12'h146B:q <= 8'h01;
            12'h146C:q <= 8'h11;
            12'h146D:q <= 8'hFF;
            12'h146E:q <= 8'h19;
            12'h146F:q <= 8'h05;
            12'h1470:q <= 8'h13;
            12'h1471:q <= 8'hFF;
            12'h1472:q <= 8'h1A;
            12'h1473:q <= 8'h1D;
            12'h1474:q <= 8'h01;
            12'h1475:q <= 8'hFF;
            12'h1476:q <= 8'h1B;
            12'h1477:q <= 8'h0F;
            12'h1478:q <= 8'h09;
            12'h1479:q <= 8'hFF;
            12'h147A:q <= 8'h1C;
            12'h147B:q <= 8'h10;
            12'h147C:q <= 8'h08;
            12'h147D:q <= 8'hFF;
            12'h147E:q <= 8'h1D;
            12'h147F:q <= 8'h1C;
            12'h1480:q <= 8'h17;
            12'h1481:q <= 8'hFF;
            12'h1482:q <= 8'h1E;
            12'h1483:q <= 8'h23;
            12'h1484:q <= 8'h19;
            12'h1485:q <= 8'hFF;
            12'h1486:q <= 8'h1F;
            12'h1487:q <= 8'h21;
            12'h1488:q <= 8'h18;
            12'h1489:q <= 8'hFF;
            12'h148A:q <= 8'h20;
            12'h148B:q <= 8'h04;
            12'h148C:q <= 8'h12;
            12'h148D:q <= 8'hFF;
            12'h148E:q <= 8'h21;
            12'h148F:q <= 8'h1E;
            12'h1490:q <= 8'h05;
            12'h1491:q <= 8'hFF;
            12'h1492:q <= 8'h22;
            12'h1493:q <= 8'h09;
            12'h1494:q <= 8'h02;
            12'h1495:q <= 8'hFF;
            12'h1496:q <= 8'h23;
            12'h1497:q <= 8'h14;
            12'h1498:q <= 8'h0F;
            12'h1499:q <= 8'hFF;
            12'h149A:q <= 8'h00;
            12'h149B:q <= 8'h0D;
            12'h149C:q <= 8'h23;
            12'h149D:q <= 8'hFF;
            12'h149E:q <= 8'h01;
            12'h149F:q <= 8'h18;
            12'h14A0:q <= 8'h1F;
            12'h14A1:q <= 8'hFF;
            12'h14A2:q <= 8'h02;
            12'h14A3:q <= 8'h1F;
            12'h14A4:q <= 8'h13;
            12'h14A5:q <= 8'hFF;
            12'h14A6:q <= 8'h03;
            12'h14A7:q <= 8'h16;
            12'h14A8:q <= 8'h0F;
            12'h14A9:q <= 8'hFF;
            12'h14AA:q <= 8'h04;
            12'h14AB:q <= 8'h08;
            12'h14AC:q <= 8'h1E;
            12'h14AD:q <= 8'hFF;
            12'h14AE:q <= 8'h05;
            12'h14AF:q <= 8'h0C;
            12'h14B0:q <= 8'h17;
            12'h14B1:q <= 8'hFF;
            12'h14B2:q <= 8'h06;
            12'h14B3:q <= 8'h1E;
            12'h14B4:q <= 8'h21;
            12'h14B5:q <= 8'hFF;
            12'h14B6:q <= 8'h07;
            12'h14B7:q <= 8'h1A;
            12'h14B8:q <= 8'h22;
            12'h14B9:q <= 8'hFF;
            12'h14BA:q <= 8'h08;
            12'h14BB:q <= 8'h07;
            12'h14BC:q <= 8'h15;
            12'h14BD:q <= 8'hFF;
            12'h14BE:q <= 8'h09;
            12'h14BF:q <= 8'h14;
            12'h14C0:q <= 8'h19;
            12'h14C1:q <= 8'hFF;
            12'h14C2:q <= 8'h0A;
            12'h14C3:q <= 8'h01;
            12'h14C4:q <= 8'h02;
            12'h14C5:q <= 8'hFF;
            12'h14C6:q <= 8'h0B;
            12'h14C7:q <= 8'h13;
            12'h14C8:q <= 8'h1A;
            12'h14C9:q <= 8'hFF;
            12'h14CA:q <= 8'h0C;
            12'h14CB:q <= 8'h1C;
            12'h14CC:q <= 8'h0A;
            12'h14CD:q <= 8'hFF;
            12'h14CE:q <= 8'h0D;
            12'h14CF:q <= 8'h0F;
            12'h14D0:q <= 8'h01;
            12'h14D1:q <= 8'hFF;
            12'h14D2:q <= 8'h0E;
            12'h14D3:q <= 8'h0A;
            12'h14D4:q <= 8'h04;
            12'h14D5:q <= 8'hFF;
            12'h14D6:q <= 8'h0F;
            12'h14D7:q <= 8'h09;
            12'h14D8:q <= 8'h12;
            12'h14D9:q <= 8'hFF;
            12'h14DA:q <= 8'h10;
            12'h14DB:q <= 8'h11;
            12'h14DC:q <= 8'h11;
            12'h14DD:q <= 8'hFF;
            12'h14DE:q <= 8'h11;
            12'h14DF:q <= 8'h02;
            12'h14E0:q <= 8'h00;
            12'h14E1:q <= 8'hFF;
            12'h14E2:q <= 8'h12;
            12'h14E3:q <= 8'h22;
            12'h14E4:q <= 8'h0B;
            12'h14E5:q <= 8'hFF;
            12'h14E6:q <= 8'h13;
            12'h14E7:q <= 8'h12;
            12'h14E8:q <= 8'h0E;
            12'h14E9:q <= 8'hFF;
            12'h14EA:q <= 8'h14;
            12'h14EB:q <= 8'h03;
            12'h14EC:q <= 8'h05;
            12'h14ED:q <= 8'hFF;
            12'h14EE:q <= 8'h15;
            12'h14EF:q <= 8'h05;
            12'h14F0:q <= 8'h03;
            12'h14F1:q <= 8'hFF;
            12'h14F2:q <= 8'h16;
            12'h14F3:q <= 8'h0E;
            12'h14F4:q <= 8'h1C;
            12'h14F5:q <= 8'hFF;
            12'h14F6:q <= 8'h17;
            12'h14F7:q <= 8'h15;
            12'h14F8:q <= 8'h0D;
            12'h14F9:q <= 8'hFF;
            12'h14FA:q <= 8'h18;
            12'h14FB:q <= 8'h06;
            12'h14FC:q <= 8'h20;
            12'h14FD:q <= 8'hFF;
            12'h14FE:q <= 8'h19;
            12'h14FF:q <= 8'h19;
            12'h1500:q <= 8'h08;
            12'h1501:q <= 8'hFF;
            12'h1502:q <= 8'h1A;
            12'h1503:q <= 8'h04;
            12'h1504:q <= 8'h0C;
            12'h1505:q <= 8'hFF;
            12'h1506:q <= 8'h1B;
            12'h1507:q <= 8'h23;
            12'h1508:q <= 8'h06;
            12'h1509:q <= 8'hFF;
            12'h150A:q <= 8'h1C;
            12'h150B:q <= 8'h0B;
            12'h150C:q <= 8'h07;
            12'h150D:q <= 8'hFF;
            12'h150E:q <= 8'h1D;
            12'h150F:q <= 8'h17;
            12'h1510:q <= 8'h18;
            12'h1511:q <= 8'hFF;
            12'h1512:q <= 8'h1E;
            12'h1513:q <= 8'h1D;
            12'h1514:q <= 8'h16;
            12'h1515:q <= 8'hFF;
            12'h1516:q <= 8'h1F;
            12'h1517:q <= 8'h00;
            12'h1518:q <= 8'h14;
            12'h1519:q <= 8'hFF;
            12'h151A:q <= 8'h20;
            12'h151B:q <= 8'h21;
            12'h151C:q <= 8'h1B;
            12'h151D:q <= 8'hFF;
            12'h151E:q <= 8'h21;
            12'h151F:q <= 8'h20;
            12'h1520:q <= 8'h10;
            12'h1521:q <= 8'hFF;
            12'h1522:q <= 8'h22;
            12'h1523:q <= 8'h1B;
            12'h1524:q <= 8'h1D;
            12'h1525:q <= 8'hFF;
            12'h1526:q <= 8'h23;
            12'h1527:q <= 8'h10;
            12'h1528:q <= 8'h09;
            12'h1529:q <= 8'hFF;
            12'h152A:q <= 8'h05;
            12'h152B:q <= 8'h06;
            12'h152C:q <= 8'h05;
            12'h152D:q <= 8'hFF;
            12'h152E:q <= 8'h06;
            12'h152F:q <= 8'h03;
            12'h1530:q <= 8'h04;
            12'h1531:q <= 8'hFF;
            12'h1532:q <= 8'h07;
            12'h1533:q <= 8'h02;
            12'h1534:q <= 8'h00;
            12'h1535:q <= 8'hFF;
            12'h1536:q <= 8'h08;
            12'h1537:q <= 8'h07;
            12'h1538:q <= 8'h09;
            12'h1539:q <= 8'hFF;
            12'h153A:q <= 8'h09;
            12'h153B:q <= 8'h08;
            12'h153C:q <= 8'h02;
            12'h153D:q <= 8'hFF;
            12'h153E:q <= 8'h00;
            12'h153F:q <= 8'h03;
            12'h1540:q <= 8'h07;
            12'h1541:q <= 8'hFF;
            12'h1542:q <= 8'h01;
            12'h1543:q <= 8'h00;
            12'h1544:q <= 8'h05;
            12'h1545:q <= 8'hFF;
            12'h1546:q <= 8'h02;
            12'h1547:q <= 8'h05;
            12'h1548:q <= 8'h04;
            12'h1549:q <= 8'hFF;
            12'h154A:q <= 8'h03;
            12'h154B:q <= 8'h09;
            12'h154C:q <= 8'h03;
            12'h154D:q <= 8'hFF;
            12'h154E:q <= 8'h04;
            12'h154F:q <= 8'h02;
            12'h1550:q <= 8'h09;
            12'h1551:q <= 8'hFF;
            12'h1552:q <= 8'h05;
            12'h1553:q <= 8'h06;
            12'h1554:q <= 8'h00;
            12'h1555:q <= 8'hFF;
            12'h1556:q <= 8'h06;
            12'h1557:q <= 8'h04;
            12'h1558:q <= 8'h06;
            12'h1559:q <= 8'hFF;
            12'h155A:q <= 8'h07;
            12'h155B:q <= 8'h01;
            12'h155C:q <= 8'h08;
            12'h155D:q <= 8'hFF;
            12'h155E:q <= 8'h08;
            12'h155F:q <= 8'h08;
            12'h1560:q <= 8'h02;
            12'h1561:q <= 8'hFF;
            12'h1562:q <= 8'h09;
            12'h1563:q <= 8'h07;
            12'h1564:q <= 8'h01;
            12'h1565:q <= 8'hFF;
            12'h1566:q <= 8'h00;
            12'h1567:q <= 8'h02;
            12'h1568:q <= 8'h07;
            12'h1569:q <= 8'hFF;
            12'h156A:q <= 8'h01;
            12'h156B:q <= 8'h00;
            12'h156C:q <= 8'h00;
            12'h156D:q <= 8'hFF;
            12'h156E:q <= 8'h02;
            12'h156F:q <= 8'h01;
            12'h1570:q <= 8'h08;
            12'h1571:q <= 8'hFF;
            12'h1572:q <= 8'h03;
            12'h1573:q <= 8'h05;
            12'h1574:q <= 8'h02;
            12'h1575:q <= 8'hFF;
            12'h1576:q <= 8'h04;
            12'h1577:q <= 8'h08;
            12'h1578:q <= 8'h09;
            12'h1579:q <= 8'hFF;
            12'h157A:q <= 8'h05;
            12'h157B:q <= 8'h03;
            12'h157C:q <= 8'h03;
            12'h157D:q <= 8'hFF;
            12'h157E:q <= 8'h06;
            12'h157F:q <= 8'h04;
            12'h1580:q <= 8'h06;
            12'h1581:q <= 8'hFF;
            12'h1582:q <= 8'h07;
            12'h1583:q <= 8'h09;
            12'h1584:q <= 8'h01;
            12'h1585:q <= 8'hFF;
            12'h1586:q <= 8'h08;
            12'h1587:q <= 8'h07;
            12'h1588:q <= 8'h04;
            12'h1589:q <= 8'hFF;
            12'h158A:q <= 8'h09;
            12'h158B:q <= 8'h06;
            12'h158C:q <= 8'h05;
            12'h158D:q <= 8'hFF;
            12'h158E:q <= 8'h00;
            12'h158F:q <= 8'h02;
            12'h1590:q <= 8'h04;
            12'h1591:q <= 8'hFF;
            12'h1592:q <= 8'h01;
            12'h1593:q <= 8'h07;
            12'h1594:q <= 8'h01;
            12'h1595:q <= 8'hFF;
            12'h1596:q <= 8'h02;
            12'h1597:q <= 8'h01;
            12'h1598:q <= 8'h00;
            12'h1599:q <= 8'hFF;
            12'h159A:q <= 8'h03;
            12'h159B:q <= 8'h03;
            12'h159C:q <= 8'h02;
            12'h159D:q <= 8'hFF;
            12'h159E:q <= 8'h04;
            12'h159F:q <= 8'h08;
            12'h15A0:q <= 8'h09;
            12'h15A1:q <= 8'hFF;
            12'h15A2:q <= 8'h05;
            12'h15A3:q <= 8'h04;
            12'h15A4:q <= 8'h03;
            12'h15A5:q <= 8'hFF;
            12'h15A6:q <= 8'h06;
            12'h15A7:q <= 8'h00;
            12'h15A8:q <= 8'h05;
            12'h15A9:q <= 8'hFF;
            12'h15AA:q <= 8'h07;
            12'h15AB:q <= 8'h09;
            12'h15AC:q <= 8'h06;
            12'h15AD:q <= 8'hFF;
            12'h15AE:q <= 8'h08;
            12'h15AF:q <= 8'h06;
            12'h15B0:q <= 8'h07;
            12'h15B1:q <= 8'hFF;
            12'h15B2:q <= 8'h09;
            12'h15B3:q <= 8'h05;
            12'h15B4:q <= 8'h08;
            12'h15B5:q <= 8'hFF;
            12'h15B6:q <= 8'h00;
            12'h15B7:q <= 8'h0C;
            12'h15B8:q <= 8'h1A;
            12'h15B9:q <= 8'h1D;
            12'h15BA:q <= 8'h10;
            12'h15BB:q <= 8'h06;
            12'h15BC:q <= 8'h16;
            12'h15BD:q <= 8'h0A;
            12'h15BE:q <= 8'h02;
            12'h15BF:q <= 8'h0F;
            12'h15C0:q <= 8'h0D;
            12'h15C1:q <= 8'h13;
            12'h15C2:q <= 8'h03;
            12'h15C3:q <= 8'hFF;
            12'h15C4:q <= 8'h01;
            12'h15C5:q <= 8'h13;
            12'h15C6:q <= 8'h10;
            12'h15C7:q <= 8'h08;
            12'h15C8:q <= 8'h0B;
            12'h15C9:q <= 8'h13;
            12'h15CA:q <= 8'h0D;
            12'h15CB:q <= 8'h07;
            12'h15CC:q <= 8'h11;
            12'h15CD:q <= 8'h1C;
            12'h15CE:q <= 8'h18;
            12'h15CF:q <= 8'h01;
            12'h15D0:q <= 8'h11;
            12'h15D1:q <= 8'hFF;
            12'h15D2:q <= 8'h02;
            12'h15D3:q <= 8'h05;
            12'h15D4:q <= 8'h09;
            12'h15D5:q <= 8'h13;
            12'h15D6:q <= 8'h01;
            12'h15D7:q <= 8'h05;
            12'h15D8:q <= 8'h07;
            12'h15D9:q <= 8'h0C;
            12'h15DA:q <= 8'h18;
            12'h15DB:q <= 8'h01;
            12'h15DC:q <= 8'h11;
            12'h15DD:q <= 8'h1D;
            12'h15DE:q <= 8'h10;
            12'h15DF:q <= 8'hFF;
            12'h15E0:q <= 8'h03;
            12'h15E1:q <= 8'h16;
            12'h15E2:q <= 8'h19;
            12'h15E3:q <= 8'h18;
            12'h15E4:q <= 8'h0A;
            12'h15E5:q <= 8'h08;
            12'h15E6:q <= 8'h12;
            12'h15E7:q <= 8'h06;
            12'h15E8:q <= 8'h19;
            12'h15E9:q <= 8'h00;
            12'h15EA:q <= 8'h07;
            12'h15EB:q <= 8'h0E;
            12'h15EC:q <= 8'h08;
            12'h15ED:q <= 8'hFF;
            12'h15EE:q <= 8'h04;
            12'h15EF:q <= 8'h09;
            12'h15F0:q <= 8'h04;
            12'h15F1:q <= 8'h05;
            12'h15F2:q <= 8'h11;
            12'h15F3:q <= 8'h03;
            12'h15F4:q <= 8'h18;
            12'h15F5:q <= 8'h1D;
            12'h15F6:q <= 8'h0D;
            12'h15F7:q <= 8'h1B;
            12'h15F8:q <= 8'h0A;
            12'h15F9:q <= 8'h1C;
            12'h15FA:q <= 8'h15;
            12'h15FB:q <= 8'hFF;
            12'h15FC:q <= 8'h05;
            12'h15FD:q <= 8'h0F;
            12'h15FE:q <= 8'h0B;
            12'h15FF:q <= 8'h12;
            12'h1600:q <= 8'h03;
            12'h1601:q <= 8'h10;
            12'h1602:q <= 8'h0F;
            12'h1603:q <= 8'h14;
            12'h1604:q <= 8'h04;
            12'h1605:q <= 8'h14;
            12'h1606:q <= 8'h0E;
            12'h1607:q <= 8'h02;
            12'h1608:q <= 8'h14;
            12'h1609:q <= 8'hFF;
            12'h160A:q <= 8'h06;
            12'h160B:q <= 8'h11;
            12'h160C:q <= 8'h15;
            12'h160D:q <= 8'h1A;
            12'h160E:q <= 8'h0E;
            12'h160F:q <= 8'h0B;
            12'h1610:q <= 8'h1D;
            12'h1611:q <= 8'h09;
            12'h1612:q <= 8'h15;
            12'h1613:q <= 8'h0B;
            12'h1614:q <= 8'h09;
            12'h1615:q <= 8'h06;
            12'h1616:q <= 8'h00;
            12'h1617:q <= 8'hFF;
            12'h1618:q <= 8'h07;
            12'h1619:q <= 8'h0D;
            12'h161A:q <= 8'h1B;
            12'h161B:q <= 8'h07;
            12'h161C:q <= 8'h0C;
            12'h161D:q <= 8'h01;
            12'h161E:q <= 8'h0E;
            12'h161F:q <= 8'h05;
            12'h1620:q <= 8'h12;
            12'h1621:q <= 8'h13;
            12'h1622:q <= 8'h06;
            12'h1623:q <= 8'h18;
            12'h1624:q <= 8'h07;
            12'h1625:q <= 8'hFF;
            12'h1626:q <= 8'h08;
            12'h1627:q <= 8'h1B;
            12'h1628:q <= 8'h05;
            12'h1629:q <= 8'h09;
            12'h162A:q <= 8'h1C;
            12'h162B:q <= 8'h14;
            12'h162C:q <= 8'h00;
            12'h162D:q <= 8'h03;
            12'h162E:q <= 8'h10;
            12'h162F:q <= 8'h15;
            12'h1630:q <= 8'h17;
            12'h1631:q <= 8'h04;
            12'h1632:q <= 8'h09;
            12'h1633:q <= 8'hFF;
            12'h1634:q <= 8'h09;
            12'h1635:q <= 8'h06;
            12'h1636:q <= 8'h0D;
            12'h1637:q <= 8'h04;
            12'h1638:q <= 8'h15;
            12'h1639:q <= 8'h11;
            12'h163A:q <= 8'h0A;
            12'h163B:q <= 8'h00;
            12'h163C:q <= 8'h0E;
            12'h163D:q <= 8'h02;
            12'h163E:q <= 8'h04;
            12'h163F:q <= 8'h16;
            12'h1640:q <= 8'h0C;
            12'h1641:q <= 8'hFF;
            12'h1642:q <= 8'h0A;
            12'h1643:q <= 8'h1C;
            12'h1644:q <= 8'h12;
            12'h1645:q <= 8'h16;
            12'h1646:q <= 8'h19;
            12'h1647:q <= 8'h17;
            12'h1648:q <= 8'h1A;
            12'h1649:q <= 8'h13;
            12'h164A:q <= 8'h1A;
            12'h164B:q <= 8'h0C;
            12'h164C:q <= 8'h1A;
            12'h164D:q <= 8'h1A;
            12'h164E:q <= 8'h0F;
            12'h164F:q <= 8'hFF;
            12'h1650:q <= 8'h0B;
            12'h1651:q <= 8'h0E;
            12'h1652:q <= 8'h03;
            12'h1653:q <= 8'h0F;
            12'h1654:q <= 8'h06;
            12'h1655:q <= 8'h0C;
            12'h1656:q <= 8'h04;
            12'h1657:q <= 8'h1C;
            12'h1658:q <= 8'h0B;
            12'h1659:q <= 8'h19;
            12'h165A:q <= 8'h1D;
            12'h165B:q <= 8'h1B;
            12'h165C:q <= 8'h12;
            12'h165D:q <= 8'hFF;
            12'h165E:q <= 8'h0C;
            12'h165F:q <= 8'h19;
            12'h1660:q <= 8'h0E;
            12'h1661:q <= 8'h0D;
            12'h1662:q <= 8'h02;
            12'h1663:q <= 8'h1B;
            12'h1664:q <= 8'h02;
            12'h1665:q <= 8'h1B;
            12'h1666:q <= 8'h08;
            12'h1667:q <= 8'h03;
            12'h1668:q <= 8'h05;
            12'h1669:q <= 8'h0B;
            12'h166A:q <= 8'h19;
            12'h166B:q <= 8'hFF;
            12'h166C:q <= 8'h0D;
            12'h166D:q <= 8'h0B;
            12'h166E:q <= 8'h16;
            12'h166F:q <= 8'h00;
            12'h1670:q <= 8'h17;
            12'h1671:q <= 8'h19;
            12'h1672:q <= 8'h09;
            12'h1673:q <= 8'h17;
            12'h1674:q <= 8'h01;
            12'h1675:q <= 8'h08;
            12'h1676:q <= 8'h16;
            12'h1677:q <= 8'h0D;
            12'h1678:q <= 8'h05;
            12'h1679:q <= 8'hFF;
            12'h167A:q <= 8'h0E;
            12'h167B:q <= 8'h00;
            12'h167C:q <= 8'h00;
            12'h167D:q <= 8'h1B;
            12'h167E:q <= 8'h14;
            12'h167F:q <= 8'h1C;
            12'h1680:q <= 8'h15;
            12'h1681:q <= 8'h0F;
            12'h1682:q <= 8'h16;
            12'h1683:q <= 8'h10;
            12'h1684:q <= 8'h12;
            12'h1685:q <= 8'h17;
            12'h1686:q <= 8'h0A;
            12'h1687:q <= 8'hFF;
            12'h1688:q <= 8'h0F;
            12'h1689:q <= 8'h04;
            12'h168A:q <= 8'h01;
            12'h168B:q <= 8'hFF;
            12'h168C:q <= 8'h10;
            12'h168D:q <= 8'h12;
            12'h168E:q <= 8'h1D;
            12'h168F:q <= 8'hFF;
            12'h1690:q <= 8'h11;
            12'h1691:q <= 8'h03;
            12'h1692:q <= 8'h06;
            12'h1693:q <= 8'hFF;
            12'h1694:q <= 8'h12;
            12'h1695:q <= 8'h0A;
            12'h1696:q <= 8'h1C;
            12'h1697:q <= 8'hFF;
            12'h1698:q <= 8'h13;
            12'h1699:q <= 8'h01;
            12'h169A:q <= 8'h17;
            12'h169B:q <= 8'hFF;
            12'h169C:q <= 8'h14;
            12'h169D:q <= 8'h18;
            12'h169E:q <= 8'h18;
            12'h169F:q <= 8'hFF;
            12'h16A0:q <= 8'h15;
            12'h16A1:q <= 8'h17;
            12'h16A2:q <= 8'h14;
            12'h16A3:q <= 8'hFF;
            12'h16A4:q <= 8'h16;
            12'h16A5:q <= 8'h07;
            12'h16A6:q <= 8'h08;
            12'h16A7:q <= 8'hFF;
            12'h16A8:q <= 8'h17;
            12'h16A9:q <= 8'h15;
            12'h16AA:q <= 8'h13;
            12'h16AB:q <= 8'hFF;
            12'h16AC:q <= 8'h18;
            12'h16AD:q <= 8'h1D;
            12'h16AE:q <= 8'h0A;
            12'h16AF:q <= 8'hFF;
            12'h16B0:q <= 8'h19;
            12'h16B1:q <= 8'h1A;
            12'h16B2:q <= 8'h0F;
            12'h16B3:q <= 8'hFF;
            12'h16B4:q <= 8'h1A;
            12'h16B5:q <= 8'h14;
            12'h16B6:q <= 8'h11;
            12'h16B7:q <= 8'hFF;
            12'h16B8:q <= 8'h1B;
            12'h16B9:q <= 8'h02;
            12'h16BA:q <= 8'h07;
            12'h16BB:q <= 8'hFF;
            12'h16BC:q <= 8'h1C;
            12'h16BD:q <= 8'h08;
            12'h16BE:q <= 8'h02;
            12'h16BF:q <= 8'hFF;
            12'h16C0:q <= 8'h1D;
            12'h16C1:q <= 8'h10;
            12'h16C2:q <= 8'h0C;
            12'h16C3:q <= 8'hFF;
            12'h16C4:q <= 8'h00;
            12'h16C5:q <= 8'h19;
            12'h16C6:q <= 8'h14;
            12'h16C7:q <= 8'hFF;
            12'h16C8:q <= 8'h01;
            12'h16C9:q <= 8'h0F;
            12'h16CA:q <= 8'h01;
            12'h16CB:q <= 8'hFF;
            12'h16CC:q <= 8'h02;
            12'h16CD:q <= 8'h0E;
            12'h16CE:q <= 8'h16;
            12'h16CF:q <= 8'hFF;
            12'h16D0:q <= 8'h03;
            12'h16D1:q <= 8'h15;
            12'h16D2:q <= 8'h15;
            12'h16D3:q <= 8'hFF;
            12'h16D4:q <= 8'h04;
            12'h16D5:q <= 8'h0A;
            12'h16D6:q <= 8'h03;
            12'h16D7:q <= 8'hFF;
            12'h16D8:q <= 8'h05;
            12'h16D9:q <= 8'h14;
            12'h16DA:q <= 8'h1C;
            12'h16DB:q <= 8'hFF;
            12'h16DC:q <= 8'h06;
            12'h16DD:q <= 8'h10;
            12'h16DE:q <= 8'h18;
            12'h16DF:q <= 8'hFF;
            12'h16E0:q <= 8'h07;
            12'h16E1:q <= 8'h0C;
            12'h16E2:q <= 8'h06;
            12'h16E3:q <= 8'hFF;
            12'h16E4:q <= 8'h08;
            12'h16E5:q <= 8'h11;
            12'h16E6:q <= 8'h12;
            12'h16E7:q <= 8'hFF;
            12'h16E8:q <= 8'h09;
            12'h16E9:q <= 8'h04;
            12'h16EA:q <= 8'h08;
            12'h16EB:q <= 8'hFF;
            12'h16EC:q <= 8'h0A;
            12'h16ED:q <= 8'h00;
            12'h16EE:q <= 8'h11;
            12'h16EF:q <= 8'hFF;
            12'h16F0:q <= 8'h0B;
            12'h16F1:q <= 8'h12;
            12'h16F2:q <= 8'h17;
            12'h16F3:q <= 8'hFF;
            12'h16F4:q <= 8'h0C;
            12'h16F5:q <= 8'h02;
            12'h16F6:q <= 8'h0D;
            12'h16F7:q <= 8'hFF;
            12'h16F8:q <= 8'h0D;
            12'h16F9:q <= 8'h0D;
            12'h16FA:q <= 8'h10;
            12'h16FB:q <= 8'hFF;
            12'h16FC:q <= 8'h0E;
            12'h16FD:q <= 8'h1B;
            12'h16FE:q <= 8'h1D;
            12'h16FF:q <= 8'hFF;
            12'h1700:q <= 8'h0F;
            12'h1701:q <= 8'h06;
            12'h1702:q <= 8'h0B;
            12'h1703:q <= 8'hFF;
            12'h1704:q <= 8'h10;
            12'h1705:q <= 8'h01;
            12'h1706:q <= 8'h0C;
            12'h1707:q <= 8'hFF;
            12'h1708:q <= 8'h11;
            12'h1709:q <= 8'h16;
            12'h170A:q <= 8'h07;
            12'h170B:q <= 8'hFF;
            12'h170C:q <= 8'h12;
            12'h170D:q <= 8'h1C;
            12'h170E:q <= 8'h05;
            12'h170F:q <= 8'hFF;
            12'h1710:q <= 8'h13;
            12'h1711:q <= 8'h1D;
            12'h1712:q <= 8'h0A;
            12'h1713:q <= 8'hFF;
            12'h1714:q <= 8'h14;
            12'h1715:q <= 8'h1A;
            12'h1716:q <= 8'h1B;
            12'h1717:q <= 8'hFF;
            12'h1718:q <= 8'h15;
            12'h1719:q <= 8'h13;
            12'h171A:q <= 8'h0F;
            12'h171B:q <= 8'hFF;
            12'h171C:q <= 8'h16;
            12'h171D:q <= 8'h07;
            12'h171E:q <= 8'h1A;
            12'h171F:q <= 8'hFF;
            12'h1720:q <= 8'h17;
            12'h1721:q <= 8'h09;
            12'h1722:q <= 8'h19;
            12'h1723:q <= 8'hFF;
            12'h1724:q <= 8'h18;
            12'h1725:q <= 8'h17;
            12'h1726:q <= 8'h00;
            12'h1727:q <= 8'hFF;
            12'h1728:q <= 8'h19;
            12'h1729:q <= 8'h05;
            12'h172A:q <= 8'h04;
            12'h172B:q <= 8'hFF;
            12'h172C:q <= 8'h1A;
            12'h172D:q <= 8'h08;
            12'h172E:q <= 8'h02;
            12'h172F:q <= 8'hFF;
            12'h1730:q <= 8'h1B;
            12'h1731:q <= 8'h18;
            12'h1732:q <= 8'h13;
            12'h1733:q <= 8'hFF;
            12'h1734:q <= 8'h1C;
            12'h1735:q <= 8'h03;
            12'h1736:q <= 8'h09;
            12'h1737:q <= 8'hFF;
            12'h1738:q <= 8'h1D;
            12'h1739:q <= 8'h0B;
            12'h173A:q <= 8'h0E;
            12'h173B:q <= 8'hFF;
            12'h173C:q <= 8'h00;
            12'h173D:q <= 8'h18;
            12'h173E:q <= 8'h13;
            12'h173F:q <= 8'hFF;
            12'h1740:q <= 8'h01;
            12'h1741:q <= 8'h10;
            12'h1742:q <= 8'h0E;
            12'h1743:q <= 8'hFF;
            12'h1744:q <= 8'h02;
            12'h1745:q <= 8'h08;
            12'h1746:q <= 8'h07;
            12'h1747:q <= 8'hFF;
            12'h1748:q <= 8'h03;
            12'h1749:q <= 8'h05;
            12'h174A:q <= 8'h0B;
            12'h174B:q <= 8'hFF;
            12'h174C:q <= 8'h04;
            12'h174D:q <= 8'h15;
            12'h174E:q <= 8'h03;
            12'h174F:q <= 8'hFF;
            12'h1750:q <= 8'h05;
            12'h1751:q <= 8'h14;
            12'h1752:q <= 8'h02;
            12'h1753:q <= 8'hFF;
            12'h1754:q <= 8'h06;
            12'h1755:q <= 8'h13;
            12'h1756:q <= 8'h1D;
            12'h1757:q <= 8'hFF;
            12'h1758:q <= 8'h07;
            12'h1759:q <= 8'h12;
            12'h175A:q <= 8'h01;
            12'h175B:q <= 8'hFF;
            12'h175C:q <= 8'h08;
            12'h175D:q <= 8'h19;
            12'h175E:q <= 8'h18;
            12'h175F:q <= 8'hFF;
            12'h1760:q <= 8'h09;
            12'h1761:q <= 8'h01;
            12'h1762:q <= 8'h11;
            12'h1763:q <= 8'hFF;
            12'h1764:q <= 8'h0A;
            12'h1765:q <= 8'h02;
            12'h1766:q <= 8'h15;
            12'h1767:q <= 8'hFF;
            12'h1768:q <= 8'h0B;
            12'h1769:q <= 8'h0E;
            12'h176A:q <= 8'h08;
            12'h176B:q <= 8'hFF;
            12'h176C:q <= 8'h0C;
            12'h176D:q <= 8'h00;
            12'h176E:q <= 8'h0F;
            12'h176F:q <= 8'hFF;
            12'h1770:q <= 8'h0D;
            12'h1771:q <= 8'h06;
            12'h1772:q <= 8'h14;
            12'h1773:q <= 8'hFF;
            12'h1774:q <= 8'h0E;
            12'h1775:q <= 8'h11;
            12'h1776:q <= 8'h1C;
            12'h1777:q <= 8'hFF;
            12'h1778:q <= 8'h0F;
            12'h1779:q <= 8'h1B;
            12'h177A:q <= 8'h19;
            12'h177B:q <= 8'hFF;
            12'h177C:q <= 8'h10;
            12'h177D:q <= 8'h0A;
            12'h177E:q <= 8'h1A;
            12'h177F:q <= 8'hFF;
            12'h1780:q <= 8'h11;
            12'h1781:q <= 8'h04;
            12'h1782:q <= 8'h09;
            12'h1783:q <= 8'hFF;
            12'h1784:q <= 8'h12;
            12'h1785:q <= 8'h1A;
            12'h1786:q <= 8'h00;
            12'h1787:q <= 8'hFF;
            12'h1788:q <= 8'h13;
            12'h1789:q <= 8'h03;
            12'h178A:q <= 8'h17;
            12'h178B:q <= 8'hFF;
            12'h178C:q <= 8'h14;
            12'h178D:q <= 8'h0F;
            12'h178E:q <= 8'h12;
            12'h178F:q <= 8'hFF;
            12'h1790:q <= 8'h15;
            12'h1791:q <= 8'h16;
            12'h1792:q <= 8'h0C;
            12'h1793:q <= 8'hFF;
            12'h1794:q <= 8'h16;
            12'h1795:q <= 8'h09;
            12'h1796:q <= 8'h10;
            12'h1797:q <= 8'hFF;
            12'h1798:q <= 8'h17;
            12'h1799:q <= 8'h07;
            12'h179A:q <= 8'h0A;
            12'h179B:q <= 8'hFF;
            12'h179C:q <= 8'h18;
            12'h179D:q <= 8'h17;
            12'h179E:q <= 8'h1B;
            12'h179F:q <= 8'hFF;
            12'h17A0:q <= 8'h19;
            12'h17A1:q <= 8'h1C;
            12'h17A2:q <= 8'h16;
            12'h17A3:q <= 8'hFF;
            12'h17A4:q <= 8'h1A;
            12'h17A5:q <= 8'h0C;
            12'h17A6:q <= 8'h06;
            12'h17A7:q <= 8'hFF;
            12'h17A8:q <= 8'h1B;
            12'h17A9:q <= 8'h0D;
            12'h17AA:q <= 8'h04;
            12'h17AB:q <= 8'hFF;
            12'h17AC:q <= 8'h1C;
            12'h17AD:q <= 8'h1D;
            12'h17AE:q <= 8'h0D;
            12'h17AF:q <= 8'hFF;
            12'h17B0:q <= 8'h1D;
            12'h17B1:q <= 8'h0B;
            12'h17B2:q <= 8'h05;
            12'h17B3:q <= 8'hFF;
            12'h17B4:q <= 8'h00;
            12'h17B5:q <= 8'h0B;
            12'h17B6:q <= 8'h03;
            12'h17B7:q <= 8'hFF;
            12'h17B8:q <= 8'h01;
            12'h17B9:q <= 8'h02;
            12'h17BA:q <= 8'h05;
            12'h17BB:q <= 8'hFF;
            12'h17BC:q <= 8'h02;
            12'h17BD:q <= 8'h1C;
            12'h17BE:q <= 8'h07;
            12'h17BF:q <= 8'hFF;
            12'h17C0:q <= 8'h03;
            12'h17C1:q <= 8'h1D;
            12'h17C2:q <= 8'h1D;
            12'h17C3:q <= 8'hFF;
            12'h17C4:q <= 8'h04;
            12'h17C5:q <= 8'h13;
            12'h17C6:q <= 8'h08;
            12'h17C7:q <= 8'hFF;
            12'h17C8:q <= 8'h05;
            12'h17C9:q <= 8'h11;
            12'h17CA:q <= 8'h1A;
            12'h17CB:q <= 8'hFF;
            12'h17CC:q <= 8'h06;
            12'h17CD:q <= 8'h18;
            12'h17CE:q <= 8'h18;
            12'h17CF:q <= 8'hFF;
            12'h17D0:q <= 8'h07;
            12'h17D1:q <= 8'h1A;
            12'h17D2:q <= 8'h00;
            12'h17D3:q <= 8'hFF;
            12'h17D4:q <= 8'h08;
            12'h17D5:q <= 8'h0C;
            12'h17D6:q <= 8'h09;
            12'h17D7:q <= 8'hFF;
            12'h17D8:q <= 8'h09;
            12'h17D9:q <= 8'h14;
            12'h17DA:q <= 8'h11;
            12'h17DB:q <= 8'hFF;
            12'h17DC:q <= 8'h0A;
            12'h17DD:q <= 8'h08;
            12'h17DE:q <= 8'h01;
            12'h17DF:q <= 8'hFF;
            12'h17E0:q <= 8'h0B;
            12'h17E1:q <= 8'h01;
            12'h17E2:q <= 8'h16;
            12'h17E3:q <= 8'hFF;
            12'h17E4:q <= 8'h0C;
            12'h17E5:q <= 8'h0D;
            12'h17E6:q <= 8'h0C;
            12'h17E7:q <= 8'hFF;
            12'h17E8:q <= 8'h0D;
            12'h17E9:q <= 8'h0A;
            12'h17EA:q <= 8'h15;
            12'h17EB:q <= 8'hFF;
            12'h17EC:q <= 8'h0E;
            12'h17ED:q <= 8'h1B;
            12'h17EE:q <= 8'h14;
            12'h17EF:q <= 8'hFF;
            12'h17F0:q <= 8'h0F;
            12'h17F1:q <= 8'h09;
            12'h17F2:q <= 8'h12;
            12'h17F3:q <= 8'hFF;
            12'h17F4:q <= 8'h10;
            12'h17F5:q <= 8'h0F;
            12'h17F6:q <= 8'h13;
            12'h17F7:q <= 8'hFF;
            12'h17F8:q <= 8'h11;
            12'h17F9:q <= 8'h06;
            12'h17FA:q <= 8'h1B;
            12'h17FB:q <= 8'hFF;
            12'h17FC:q <= 8'h12;
            12'h17FD:q <= 8'h10;
            12'h17FE:q <= 8'h0F;
            12'h17FF:q <= 8'hFF;
            12'h1800:q <= 8'h13;
            12'h1801:q <= 8'h16;
            12'h1802:q <= 8'h04;
            12'h1803:q <= 8'hFF;
            12'h1804:q <= 8'h14;
            12'h1805:q <= 8'h19;
            12'h1806:q <= 8'h1C;
            12'h1807:q <= 8'hFF;
            12'h1808:q <= 8'h15;
            12'h1809:q <= 8'h03;
            12'h180A:q <= 8'h06;
            12'h180B:q <= 8'hFF;
            12'h180C:q <= 8'h16;
            12'h180D:q <= 8'h15;
            12'h180E:q <= 8'h17;
            12'h180F:q <= 8'hFF;
            12'h1810:q <= 8'h17;
            12'h1811:q <= 8'h04;
            12'h1812:q <= 8'h0E;
            12'h1813:q <= 8'hFF;
            12'h1814:q <= 8'h18;
            12'h1815:q <= 8'h17;
            12'h1816:q <= 8'h10;
            12'h1817:q <= 8'hFF;
            12'h1818:q <= 8'h19;
            12'h1819:q <= 8'h05;
            12'h181A:q <= 8'h0B;
            12'h181B:q <= 8'hFF;
            12'h181C:q <= 8'h1A;
            12'h181D:q <= 8'h07;
            12'h181E:q <= 8'h02;
            12'h181F:q <= 8'hFF;
            12'h1820:q <= 8'h1B;
            12'h1821:q <= 8'h0E;
            12'h1822:q <= 8'h0A;
            12'h1823:q <= 8'hFF;
            12'h1824:q <= 8'h1C;
            12'h1825:q <= 8'h00;
            12'h1826:q <= 8'h19;
            12'h1827:q <= 8'hFF;
            12'h1828:q <= 8'h1D;
            12'h1829:q <= 8'h12;
            12'h182A:q <= 8'h0D;
            12'h182B:q <= 8'hFF;
            12'h182C:q <= 8'h00;
            12'h182D:q <= 8'h1D;
            12'h182E:q <= 8'h07;
            12'h182F:q <= 8'hFF;
            12'h1830:q <= 8'h01;
            12'h1831:q <= 8'h15;
            12'h1832:q <= 8'h09;
            12'h1833:q <= 8'hFF;
            12'h1834:q <= 8'h02;
            12'h1835:q <= 8'h14;
            12'h1836:q <= 8'h13;
            12'h1837:q <= 8'hFF;
            12'h1838:q <= 8'h03;
            12'h1839:q <= 8'h07;
            12'h183A:q <= 8'h12;
            12'h183B:q <= 8'hFF;
            12'h183C:q <= 8'h04;
            12'h183D:q <= 8'h18;
            12'h183E:q <= 8'h14;
            12'h183F:q <= 8'hFF;
            12'h1840:q <= 8'h05;
            12'h1841:q <= 8'h0E;
            12'h1842:q <= 8'h1D;
            12'h1843:q <= 8'hFF;
            12'h1844:q <= 8'h06;
            12'h1845:q <= 8'h0F;
            12'h1846:q <= 8'h15;
            12'h1847:q <= 8'hFF;
            12'h1848:q <= 8'h07;
            12'h1849:q <= 8'h1C;
            12'h184A:q <= 8'h0E;
            12'h184B:q <= 8'hFF;
            12'h184C:q <= 8'h08;
            12'h184D:q <= 8'h0A;
            12'h184E:q <= 8'h1C;
            12'h184F:q <= 8'hFF;
            12'h1850:q <= 8'h09;
            12'h1851:q <= 8'h10;
            12'h1852:q <= 8'h06;
            12'h1853:q <= 8'hFF;
            12'h1854:q <= 8'h0A;
            12'h1855:q <= 8'h08;
            12'h1856:q <= 8'h02;
            12'h1857:q <= 8'hFF;
            12'h1858:q <= 8'h0B;
            12'h1859:q <= 8'h01;
            12'h185A:q <= 8'h1B;
            12'h185B:q <= 8'hFF;
            12'h185C:q <= 8'h0C;
            12'h185D:q <= 8'h02;
            12'h185E:q <= 8'h05;
            12'h185F:q <= 8'hFF;
            12'h1860:q <= 8'h0D;
            12'h1861:q <= 8'h09;
            12'h1862:q <= 8'h0A;
            12'h1863:q <= 8'hFF;
            12'h1864:q <= 8'h0E;
            12'h1865:q <= 8'h12;
            12'h1866:q <= 8'h16;
            12'h1867:q <= 8'hFF;
            12'h1868:q <= 8'h0F;
            12'h1869:q <= 8'h17;
            12'h186A:q <= 8'h0C;
            12'h186B:q <= 8'hFF;
            12'h186C:q <= 8'h10;
            12'h186D:q <= 8'h00;
            12'h186E:q <= 8'h0F;
            12'h186F:q <= 8'hFF;
            12'h1870:q <= 8'h11;
            12'h1871:q <= 8'h04;
            12'h1872:q <= 8'h03;
            12'h1873:q <= 8'hFF;
            12'h1874:q <= 8'h12;
            12'h1875:q <= 8'h1A;
            12'h1876:q <= 8'h10;
            12'h1877:q <= 8'hFF;
            12'h1878:q <= 8'h13;
            12'h1879:q <= 8'h11;
            12'h187A:q <= 8'h19;
            12'h187B:q <= 8'hFF;
            12'h187C:q <= 8'h14;
            12'h187D:q <= 8'h13;
            12'h187E:q <= 8'h00;
            12'h187F:q <= 8'hFF;
            12'h1880:q <= 8'h15;
            12'h1881:q <= 8'h16;
            12'h1882:q <= 8'h08;
            12'h1883:q <= 8'hFF;
            12'h1884:q <= 8'h16;
            12'h1885:q <= 8'h0D;
            12'h1886:q <= 8'h18;
            12'h1887:q <= 8'hFF;
            12'h1888:q <= 8'h17;
            12'h1889:q <= 8'h06;
            12'h188A:q <= 8'h17;
            12'h188B:q <= 8'hFF;
            12'h188C:q <= 8'h18;
            12'h188D:q <= 8'h0B;
            12'h188E:q <= 8'h0D;
            12'h188F:q <= 8'hFF;
            12'h1890:q <= 8'h19;
            12'h1891:q <= 8'h19;
            12'h1892:q <= 8'h0B;
            12'h1893:q <= 8'hFF;
            12'h1894:q <= 8'h1A;
            12'h1895:q <= 8'h0C;
            12'h1896:q <= 8'h04;
            12'h1897:q <= 8'hFF;
            12'h1898:q <= 8'h1B;
            12'h1899:q <= 8'h05;
            12'h189A:q <= 8'h1A;
            12'h189B:q <= 8'hFF;
            12'h189C:q <= 8'h1C;
            12'h189D:q <= 8'h03;
            12'h189E:q <= 8'h01;
            12'h189F:q <= 8'hFF;
            12'h18A0:q <= 8'h1D;
            12'h18A1:q <= 8'h1B;
            12'h18A2:q <= 8'h11;
            12'h18A3:q <= 8'hFF;
            12'h18A4:q <= 8'h03;
            12'h18A5:q <= 8'h01;
            12'h18A6:q <= 8'h03;
            12'h18A7:q <= 8'h01;
            12'h18A8:q <= 8'h04;
            12'h18A9:q <= 8'h07;
            12'h18AA:q <= 8'h04;
            12'h18AB:q <= 8'h06;
            12'h18AC:q <= 8'h05;
            12'h18AD:q <= 8'h04;
            12'h18AE:q <= 8'h00;
            12'h18AF:q <= 8'h06;
            12'h18B0:q <= 8'h05;
            12'h18B1:q <= 8'hFF;
            12'h18B2:q <= 8'h04;
            12'h18B3:q <= 8'h07;
            12'h18B4:q <= 8'h06;
            12'h18B5:q <= 8'hFF;
            12'h18B6:q <= 8'h05;
            12'h18B7:q <= 8'h06;
            12'h18B8:q <= 8'h00;
            12'h18B9:q <= 8'hFF;
            12'h18BA:q <= 8'h06;
            12'h18BB:q <= 8'h02;
            12'h18BC:q <= 8'h02;
            12'h18BD:q <= 8'hFF;
            12'h18BE:q <= 8'h07;
            12'h18BF:q <= 8'h04;
            12'h18C0:q <= 8'h05;
            12'h18C1:q <= 8'hFF;
            12'h18C2:q <= 8'h00;
            12'h18C3:q <= 8'h07;
            12'h18C4:q <= 8'h00;
            12'h18C5:q <= 8'hFF;
            12'h18C6:q <= 8'h01;
            12'h18C7:q <= 8'h06;
            12'h18C8:q <= 8'h04;
            12'h18C9:q <= 8'hFF;
            12'h18CA:q <= 8'h02;
            12'h18CB:q <= 8'h01;
            12'h18CC:q <= 8'h03;
            12'h18CD:q <= 8'hFF;
            12'h18CE:q <= 8'h03;
            12'h18CF:q <= 8'h00;
            12'h18D0:q <= 8'h07;
            12'h18D1:q <= 8'hFF;
            12'h18D2:q <= 8'h04;
            12'h18D3:q <= 8'h05;
            12'h18D4:q <= 8'h02;
            12'h18D5:q <= 8'hFF;
            12'h18D6:q <= 8'h05;
            12'h18D7:q <= 8'h04;
            12'h18D8:q <= 8'h06;
            12'h18D9:q <= 8'hFF;
            12'h18DA:q <= 8'h06;
            12'h18DB:q <= 8'h02;
            12'h18DC:q <= 8'h05;
            12'h18DD:q <= 8'hFF;
            12'h18DE:q <= 8'h07;
            12'h18DF:q <= 8'h03;
            12'h18E0:q <= 8'h01;
            12'h18E1:q <= 8'hFF;
            12'h18E2:q <= 8'h00;
            12'h18E3:q <= 8'h05;
            12'h18E4:q <= 8'h05;
            12'h18E5:q <= 8'hFF;
            12'h18E6:q <= 8'h01;
            12'h18E7:q <= 8'h07;
            12'h18E8:q <= 8'h01;
            12'h18E9:q <= 8'hFF;
            12'h18EA:q <= 8'h02;
            12'h18EB:q <= 8'h00;
            12'h18EC:q <= 8'h00;
            12'h18ED:q <= 8'hFF;
            12'h18EE:q <= 8'h03;
            12'h18EF:q <= 8'h02;
            12'h18F0:q <= 8'h07;
            12'h18F1:q <= 8'hFF;
            12'h18F2:q <= 8'h04;
            12'h18F3:q <= 8'h04;
            12'h18F4:q <= 8'h02;
            12'h18F5:q <= 8'hFF;
            12'h18F6:q <= 8'h05;
            12'h18F7:q <= 8'h03;
            12'h18F8:q <= 8'h06;
            12'h18F9:q <= 8'hFF;
            12'h18FA:q <= 8'h06;
            12'h18FB:q <= 8'h01;
            12'h18FC:q <= 8'h04;
            12'h18FD:q <= 8'hFF;
            12'h18FE:q <= 8'h07;
            12'h18FF:q <= 8'h06;
            12'h1900:q <= 8'h03;
            12'h1901:q <= 8'hFF;
            12'h1902:q <= 8'h00;
            12'h1903:q <= 8'h02;
            12'h1904:q <= 8'h00;
            12'h1905:q <= 8'hFF;
            12'h1906:q <= 8'h01;
            12'h1907:q <= 8'h05;
            12'h1908:q <= 8'h05;
            12'h1909:q <= 8'hFF;
            12'h190A:q <= 8'h02;
            12'h190B:q <= 8'h01;
            12'h190C:q <= 8'h02;
            12'h190D:q <= 8'hFF;
            12'h190E:q <= 8'h03;
            12'h190F:q <= 8'h06;
            12'h1910:q <= 8'h01;
            12'h1911:q <= 8'hFF;
            12'h1912:q <= 8'h04;
            12'h1913:q <= 8'h07;
            12'h1914:q <= 8'h04;
            12'h1915:q <= 8'hFF;
            12'h1916:q <= 8'h05;
            12'h1917:q <= 8'h00;
            12'h1918:q <= 8'h03;
            12'h1919:q <= 8'hFF;
            12'h191A:q <= 8'h06;
            12'h191B:q <= 8'h03;
            12'h191C:q <= 8'h06;
            12'h191D:q <= 8'hFF;
            12'h191E:q <= 8'h07;
            12'h191F:q <= 8'h04;
            12'h1920:q <= 8'h07;
            12'h1921:q <= 8'hFF;
            12'h1922:q <= 8'h00;
            12'h1923:q <= 8'h05;
            12'h1924:q <= 8'h01;
            12'h1925:q <= 8'hFF;
            12'h1926:q <= 8'h01;
            12'h1927:q <= 8'h01;
            12'h1928:q <= 8'h03;
            12'h1929:q <= 8'hFF;
            12'h192A:q <= 8'h02;
            12'h192B:q <= 8'h06;
            12'h192C:q <= 8'h02;
            12'h192D:q <= 8'hFF;
            12'h192E:q <= 8'h03;
            12'h192F:q <= 8'h07;
            12'h1930:q <= 8'h06;
            12'h1931:q <= 8'hFF;
            12'h1932:q <= 8'h04;
            12'h1933:q <= 8'h02;
            12'h1934:q <= 8'h04;
            12'h1935:q <= 8'hFF;
            12'h1936:q <= 8'h05;
            12'h1937:q <= 8'h00;
            12'h1938:q <= 8'h07;
            12'h1939:q <= 8'hFF;
            12'h193A:q <= 8'h06;
            12'h193B:q <= 8'h03;
            12'h193C:q <= 8'h05;
            12'h193D:q <= 8'hFF;
            12'h193E:q <= 8'h07;
            12'h193F:q <= 8'h04;
            12'h1940:q <= 8'h00;
            12'h1941:q <= 8'hFF;
            12'h1942:q <= 8'h00;
            12'h1943:q <= 8'h0F;
            12'h1944:q <= 8'h08;
            12'h1945:q <= 8'h02;
            12'h1946:q <= 8'hFF;
            12'h1947:q <= 8'h01;
            12'h1948:q <= 8'h00;
            12'h1949:q <= 8'h0C;
            12'h194A:q <= 8'h08;
            12'h194B:q <= 8'hFF;
            12'h194C:q <= 8'h02;
            12'h194D:q <= 8'h11;
            12'h194E:q <= 8'h07;
            12'h194F:q <= 8'h0A;
            12'h1950:q <= 8'hFF;
            12'h1951:q <= 8'h03;
            12'h1952:q <= 8'h01;
            12'h1953:q <= 8'h10;
            12'h1954:q <= 8'h13;
            12'h1955:q <= 8'hFF;
            12'h1956:q <= 8'h04;
            12'h1957:q <= 8'h0C;
            12'h1958:q <= 8'h11;
            12'h1959:q <= 8'h04;
            12'h195A:q <= 8'hFF;
            12'h195B:q <= 8'h05;
            12'h195C:q <= 8'h07;
            12'h195D:q <= 8'h05;
            12'h195E:q <= 8'h03;
            12'h195F:q <= 8'hFF;
            12'h1960:q <= 8'h06;
            12'h1961:q <= 8'h0E;
            12'h1962:q <= 8'h09;
            12'h1963:q <= 8'h0F;
            12'h1964:q <= 8'hFF;
            12'h1965:q <= 8'h07;
            12'h1966:q <= 8'h0A;
            12'h1967:q <= 8'h02;
            12'h1968:q <= 8'h0E;
            12'h1969:q <= 8'hFF;
            12'h196A:q <= 8'h08;
            12'h196B:q <= 8'h08;
            12'h196C:q <= 8'h0D;
            12'h196D:q <= 8'h01;
            12'h196E:q <= 8'hFF;
            12'h196F:q <= 8'h09;
            12'h1970:q <= 8'h06;
            12'h1971:q <= 8'h04;
            12'h1972:q <= 8'h07;
            12'h1973:q <= 8'hFF;
            12'h1974:q <= 8'h0A;
            12'h1975:q <= 8'h10;
            12'h1976:q <= 8'h0A;
            12'h1977:q <= 8'h0D;
            12'h1978:q <= 8'hFF;
            12'h1979:q <= 8'h0B;
            12'h197A:q <= 8'h0D;
            12'h197B:q <= 8'h13;
            12'h197C:q <= 8'h0B;
            12'h197D:q <= 8'hFF;
            12'h197E:q <= 8'h0C;
            12'h197F:q <= 8'h05;
            12'h1980:q <= 8'h06;
            12'h1981:q <= 8'h05;
            12'h1982:q <= 8'hFF;
            12'h1983:q <= 8'h0D;
            12'h1984:q <= 8'h03;
            12'h1985:q <= 8'h03;
            12'h1986:q <= 8'h09;
            12'h1987:q <= 8'hFF;
            12'h1988:q <= 8'h0E;
            12'h1989:q <= 8'h09;
            12'h198A:q <= 8'h0F;
            12'h198B:q <= 8'h0C;
            12'h198C:q <= 8'hFF;
            12'h198D:q <= 8'h0F;
            12'h198E:q <= 8'h13;
            12'h198F:q <= 8'h00;
            12'h1990:q <= 8'h11;
            12'h1991:q <= 8'hFF;
            12'h1992:q <= 8'h10;
            12'h1993:q <= 8'h04;
            12'h1994:q <= 8'h0B;
            12'h1995:q <= 8'h12;
            12'h1996:q <= 8'hFF;
            12'h1997:q <= 8'h11;
            12'h1998:q <= 8'h02;
            12'h1999:q <= 8'h01;
            12'h199A:q <= 8'h00;
            12'h199B:q <= 8'hFF;
            12'h199C:q <= 8'h12;
            12'h199D:q <= 8'h0B;
            12'h199E:q <= 8'h0E;
            12'h199F:q <= 8'h10;
            12'h19A0:q <= 8'hFF;
            12'h19A1:q <= 8'h13;
            12'h19A2:q <= 8'h12;
            12'h19A3:q <= 8'h12;
            12'h19A4:q <= 8'h06;
            12'h19A5:q <= 8'hFF;
            12'h19A6:q <= 8'h00;
            12'h19A7:q <= 8'h10;
            12'h19A8:q <= 8'h06;
            12'h19A9:q <= 8'hFF;
            12'h19AA:q <= 8'h01;
            12'h19AB:q <= 8'h04;
            12'h19AC:q <= 8'h10;
            12'h19AD:q <= 8'hFF;
            12'h19AE:q <= 8'h02;
            12'h19AF:q <= 8'h0A;
            12'h19B0:q <= 8'h04;
            12'h19B1:q <= 8'hFF;
            12'h19B2:q <= 8'h03;
            12'h19B3:q <= 8'h07;
            12'h19B4:q <= 8'h07;
            12'h19B5:q <= 8'hFF;
            12'h19B6:q <= 8'h04;
            12'h19B7:q <= 8'h12;
            12'h19B8:q <= 8'h13;
            12'h19B9:q <= 8'hFF;
            12'h19BA:q <= 8'h05;
            12'h19BB:q <= 8'h00;
            12'h19BC:q <= 8'h0A;
            12'h19BD:q <= 8'hFF;
            12'h19BE:q <= 8'h06;
            12'h19BF:q <= 8'h03;
            12'h19C0:q <= 8'h0B;
            12'h19C1:q <= 8'hFF;
            12'h19C2:q <= 8'h07;
            12'h19C3:q <= 8'h13;
            12'h19C4:q <= 8'h05;
            12'h19C5:q <= 8'hFF;
            12'h19C6:q <= 8'h08;
            12'h19C7:q <= 8'h11;
            12'h19C8:q <= 8'h0D;
            12'h19C9:q <= 8'hFF;
            12'h19CA:q <= 8'h09;
            12'h19CB:q <= 8'h08;
            12'h19CC:q <= 8'h02;
            12'h19CD:q <= 8'hFF;
            12'h19CE:q <= 8'h0A;
            12'h19CF:q <= 8'h01;
            12'h19D0:q <= 8'h0F;
            12'h19D1:q <= 8'hFF;
            12'h19D2:q <= 8'h0B;
            12'h19D3:q <= 8'h05;
            12'h19D4:q <= 8'h0E;
            12'h19D5:q <= 8'hFF;
            12'h19D6:q <= 8'h0C;
            12'h19D7:q <= 8'h06;
            12'h19D8:q <= 8'h0C;
            12'h19D9:q <= 8'hFF;
            12'h19DA:q <= 8'h0D;
            12'h19DB:q <= 8'h09;
            12'h19DC:q <= 8'h09;
            12'h19DD:q <= 8'hFF;
            12'h19DE:q <= 8'h0E;
            12'h19DF:q <= 8'h0B;
            12'h19E0:q <= 8'h00;
            12'h19E1:q <= 8'hFF;
            12'h19E2:q <= 8'h0F;
            12'h19E3:q <= 8'h0C;
            12'h19E4:q <= 8'h01;
            12'h19E5:q <= 8'hFF;
            12'h19E6:q <= 8'h10;
            12'h19E7:q <= 8'h0F;
            12'h19E8:q <= 8'h03;
            12'h19E9:q <= 8'hFF;
            12'h19EA:q <= 8'h11;
            12'h19EB:q <= 8'h0D;
            12'h19EC:q <= 8'h11;
            12'h19ED:q <= 8'hFF;
            12'h19EE:q <= 8'h12;
            12'h19EF:q <= 8'h02;
            12'h19F0:q <= 8'h12;
            12'h19F1:q <= 8'hFF;
            12'h19F2:q <= 8'h13;
            12'h19F3:q <= 8'h0E;
            12'h19F4:q <= 8'h08;
            12'h19F5:q <= 8'hFF;
            12'h19F6:q <= 8'h00;
            12'h19F7:q <= 8'h10;
            12'h19F8:q <= 8'h06;
            12'h19F9:q <= 8'hFF;
            12'h19FA:q <= 8'h01;
            12'h19FB:q <= 8'h0D;
            12'h19FC:q <= 8'h09;
            12'h19FD:q <= 8'hFF;
            12'h19FE:q <= 8'h02;
            12'h19FF:q <= 8'h0A;
            12'h1A00:q <= 8'h0E;
            12'h1A01:q <= 8'hFF;
            12'h1A02:q <= 8'h03;
            12'h1A03:q <= 8'h02;
            12'h1A04:q <= 8'h01;
            12'h1A05:q <= 8'hFF;
            12'h1A06:q <= 8'h04;
            12'h1A07:q <= 8'h05;
            12'h1A08:q <= 8'h04;
            12'h1A09:q <= 8'hFF;
            12'h1A0A:q <= 8'h05;
            12'h1A0B:q <= 8'h0B;
            12'h1A0C:q <= 8'h03;
            12'h1A0D:q <= 8'hFF;
            12'h1A0E:q <= 8'h06;
            12'h1A0F:q <= 8'h0C;
            12'h1A10:q <= 8'h0C;
            12'h1A11:q <= 8'hFF;
            12'h1A12:q <= 8'h07;
            12'h1A13:q <= 8'h0F;
            12'h1A14:q <= 8'h0F;
            12'h1A15:q <= 8'hFF;
            12'h1A16:q <= 8'h08;
            12'h1A17:q <= 8'h11;
            12'h1A18:q <= 8'h0B;
            12'h1A19:q <= 8'hFF;
            12'h1A1A:q <= 8'h09;
            12'h1A1B:q <= 8'h06;
            12'h1A1C:q <= 8'h0A;
            12'h1A1D:q <= 8'hFF;
            12'h1A1E:q <= 8'h0A;
            12'h1A1F:q <= 8'h09;
            12'h1A20:q <= 8'h00;
            12'h1A21:q <= 8'hFF;
            12'h1A22:q <= 8'h0B;
            12'h1A23:q <= 8'h04;
            12'h1A24:q <= 8'h08;
            12'h1A25:q <= 8'hFF;
            12'h1A26:q <= 8'h0C;
            12'h1A27:q <= 8'h08;
            12'h1A28:q <= 8'h13;
            12'h1A29:q <= 8'hFF;
            12'h1A2A:q <= 8'h0D;
            12'h1A2B:q <= 8'h03;
            12'h1A2C:q <= 8'h10;
            12'h1A2D:q <= 8'hFF;
            12'h1A2E:q <= 8'h0E;
            12'h1A2F:q <= 8'h07;
            12'h1A30:q <= 8'h0D;
            12'h1A31:q <= 8'hFF;
            12'h1A32:q <= 8'h0F;
            12'h1A33:q <= 8'h0E;
            12'h1A34:q <= 8'h02;
            12'h1A35:q <= 8'hFF;
            12'h1A36:q <= 8'h10;
            12'h1A37:q <= 8'h12;
            12'h1A38:q <= 8'h05;
            12'h1A39:q <= 8'hFF;
            12'h1A3A:q <= 8'h11;
            12'h1A3B:q <= 8'h00;
            12'h1A3C:q <= 8'h11;
            12'h1A3D:q <= 8'hFF;
            12'h1A3E:q <= 8'h12;
            12'h1A3F:q <= 8'h13;
            12'h1A40:q <= 8'h12;
            12'h1A41:q <= 8'hFF;
            12'h1A42:q <= 8'h13;
            12'h1A43:q <= 8'h01;
            12'h1A44:q <= 8'h07;
            12'h1A45:q <= 8'hFF;
            12'h1A46:q <= 8'h00;
            12'h1A47:q <= 8'h08;
            12'h1A48:q <= 8'h06;
            12'h1A49:q <= 8'hFF;
            12'h1A4A:q <= 8'h01;
            12'h1A4B:q <= 8'h06;
            12'h1A4C:q <= 8'h05;
            12'h1A4D:q <= 8'hFF;
            12'h1A4E:q <= 8'h02;
            12'h1A4F:q <= 8'h13;
            12'h1A50:q <= 8'h0B;
            12'h1A51:q <= 8'hFF;
            12'h1A52:q <= 8'h03;
            12'h1A53:q <= 8'h03;
            12'h1A54:q <= 8'h01;
            12'h1A55:q <= 8'hFF;
            12'h1A56:q <= 8'h04;
            12'h1A57:q <= 8'h0E;
            12'h1A58:q <= 8'h07;
            12'h1A59:q <= 8'hFF;
            12'h1A5A:q <= 8'h05;
            12'h1A5B:q <= 8'h11;
            12'h1A5C:q <= 8'h13;
            12'h1A5D:q <= 8'hFF;
            12'h1A5E:q <= 8'h06;
            12'h1A5F:q <= 8'h01;
            12'h1A60:q <= 8'h0C;
            12'h1A61:q <= 8'hFF;
            12'h1A62:q <= 8'h07;
            12'h1A63:q <= 8'h10;
            12'h1A64:q <= 8'h10;
            12'h1A65:q <= 8'hFF;
            12'h1A66:q <= 8'h08;
            12'h1A67:q <= 8'h0A;
            12'h1A68:q <= 8'h12;
            12'h1A69:q <= 8'hFF;
            12'h1A6A:q <= 8'h09;
            12'h1A6B:q <= 8'h0B;
            12'h1A6C:q <= 8'h0E;
            12'h1A6D:q <= 8'hFF;
            12'h1A6E:q <= 8'h0A;
            12'h1A6F:q <= 8'h07;
            12'h1A70:q <= 8'h08;
            12'h1A71:q <= 8'hFF;
            12'h1A72:q <= 8'h0B;
            12'h1A73:q <= 8'h04;
            12'h1A74:q <= 8'h0F;
            12'h1A75:q <= 8'hFF;
            12'h1A76:q <= 8'h0C;
            12'h1A77:q <= 8'h02;
            12'h1A78:q <= 8'h09;
            12'h1A79:q <= 8'hFF;
            12'h1A7A:q <= 8'h0D;
            12'h1A7B:q <= 8'h0C;
            12'h1A7C:q <= 8'h0D;
            12'h1A7D:q <= 8'hFF;
            12'h1A7E:q <= 8'h0E;
            12'h1A7F:q <= 8'h0D;
            12'h1A80:q <= 8'h04;
            12'h1A81:q <= 8'hFF;
            12'h1A82:q <= 8'h0F;
            12'h1A83:q <= 8'h0F;
            12'h1A84:q <= 8'h0A;
            12'h1A85:q <= 8'hFF;
            12'h1A86:q <= 8'h10;
            12'h1A87:q <= 8'h05;
            12'h1A88:q <= 8'h02;
            12'h1A89:q <= 8'hFF;
            12'h1A8A:q <= 8'h11;
            12'h1A8B:q <= 8'h12;
            12'h1A8C:q <= 8'h00;
            12'h1A8D:q <= 8'hFF;
            12'h1A8E:q <= 8'h12;
            12'h1A8F:q <= 8'h09;
            12'h1A90:q <= 8'h11;
            12'h1A91:q <= 8'hFF;
            12'h1A92:q <= 8'h13;
            12'h1A93:q <= 8'h00;
            12'h1A94:q <= 8'h03;
            12'h1A95:q <= 8'hFF;
            12'h1A96:q <= 8'h00;
            12'h1A97:q <= 8'h09;
            12'h1A98:q <= 8'h0B;
            12'h1A99:q <= 8'hFF;
            12'h1A9A:q <= 8'h01;
            12'h1A9B:q <= 8'h11;
            12'h1A9C:q <= 8'h04;
            12'h1A9D:q <= 8'hFF;
            12'h1A9E:q <= 8'h02;
            12'h1A9F:q <= 8'h08;
            12'h1AA0:q <= 8'h03;
            12'h1AA1:q <= 8'hFF;
            12'h1AA2:q <= 8'h03;
            12'h1AA3:q <= 8'h12;
            12'h1AA4:q <= 8'h00;
            12'h1AA5:q <= 8'hFF;
            12'h1AA6:q <= 8'h04;
            12'h1AA7:q <= 8'h06;
            12'h1AA8:q <= 8'h0F;
            12'h1AA9:q <= 8'hFF;
            12'h1AAA:q <= 8'h05;
            12'h1AAB:q <= 8'h0F;
            12'h1AAC:q <= 8'h0E;
            12'h1AAD:q <= 8'hFF;
            12'h1AAE:q <= 8'h06;
            12'h1AAF:q <= 8'h01;
            12'h1AB0:q <= 8'h07;
            12'h1AB1:q <= 8'hFF;
            12'h1AB2:q <= 8'h07;
            12'h1AB3:q <= 8'h0D;
            12'h1AB4:q <= 8'h0C;
            12'h1AB5:q <= 8'hFF;
            12'h1AB6:q <= 8'h08;
            12'h1AB7:q <= 8'h07;
            12'h1AB8:q <= 8'h09;
            12'h1AB9:q <= 8'hFF;
            12'h1ABA:q <= 8'h09;
            12'h1ABB:q <= 8'h13;
            12'h1ABC:q <= 8'h05;
            12'h1ABD:q <= 8'hFF;
            12'h1ABE:q <= 8'h0A;
            12'h1ABF:q <= 8'h03;
            12'h1AC0:q <= 8'h08;
            12'h1AC1:q <= 8'hFF;
            12'h1AC2:q <= 8'h0B;
            12'h1AC3:q <= 8'h00;
            12'h1AC4:q <= 8'h02;
            12'h1AC5:q <= 8'hFF;
            12'h1AC6:q <= 8'h0C;
            12'h1AC7:q <= 8'h0E;
            12'h1AC8:q <= 8'h01;
            12'h1AC9:q <= 8'hFF;
            12'h1ACA:q <= 8'h0D;
            12'h1ACB:q <= 8'h04;
            12'h1ACC:q <= 8'h0A;
            12'h1ACD:q <= 8'hFF;
            12'h1ACE:q <= 8'h0E;
            12'h1ACF:q <= 8'h05;
            12'h1AD0:q <= 8'h0D;
            12'h1AD1:q <= 8'hFF;
            12'h1AD2:q <= 8'h0F;
            12'h1AD3:q <= 8'h0B;
            12'h1AD4:q <= 8'h06;
            12'h1AD5:q <= 8'hFF;
            12'h1AD6:q <= 8'h10;
            12'h1AD7:q <= 8'h0A;
            12'h1AD8:q <= 8'h10;
            12'h1AD9:q <= 8'hFF;
            12'h1ADA:q <= 8'h11;
            12'h1ADB:q <= 8'h0C;
            12'h1ADC:q <= 8'h12;
            12'h1ADD:q <= 8'hFF;
            12'h1ADE:q <= 8'h12;
            12'h1ADF:q <= 8'h02;
            12'h1AE0:q <= 8'h11;
            12'h1AE1:q <= 8'hFF;
            12'h1AE2:q <= 8'h13;
            12'h1AE3:q <= 8'h10;
            12'h1AE4:q <= 8'h13;
            12'h1AE5:q <= 8'hFF;
            12'h1AE6:q <= 8'h00;
            12'h1AE7:q <= 8'h0A;
            12'h1AE8:q <= 8'h0C;
            12'h1AE9:q <= 8'hFF;
            12'h1AEA:q <= 8'h01;
            12'h1AEB:q <= 8'h02;
            12'h1AEC:q <= 8'h13;
            12'h1AED:q <= 8'hFF;
            12'h1AEE:q <= 8'h02;
            12'h1AEF:q <= 8'h11;
            12'h1AF0:q <= 8'h0A;
            12'h1AF1:q <= 8'hFF;
            12'h1AF2:q <= 8'h03;
            12'h1AF3:q <= 8'h08;
            12'h1AF4:q <= 8'h0D;
            12'h1AF5:q <= 8'hFF;
            12'h1AF6:q <= 8'h04;
            12'h1AF7:q <= 8'h13;
            12'h1AF8:q <= 8'h11;
            12'h1AF9:q <= 8'hFF;
            12'h1AFA:q <= 8'h05;
            12'h1AFB:q <= 8'h10;
            12'h1AFC:q <= 8'h02;
            12'h1AFD:q <= 8'hFF;
            12'h1AFE:q <= 8'h06;
            12'h1AFF:q <= 8'h0F;
            12'h1B00:q <= 8'h06;
            12'h1B01:q <= 8'hFF;
            12'h1B02:q <= 8'h07;
            12'h1B03:q <= 8'h0B;
            12'h1B04:q <= 8'h08;
            12'h1B05:q <= 8'hFF;
            12'h1B06:q <= 8'h08;
            12'h1B07:q <= 8'h12;
            12'h1B08:q <= 8'h01;
            12'h1B09:q <= 8'hFF;
            12'h1B0A:q <= 8'h09;
            12'h1B0B:q <= 8'h00;
            12'h1B0C:q <= 8'h00;
            12'h1B0D:q <= 8'hFF;
            12'h1B0E:q <= 8'h0A;
            12'h1B0F:q <= 8'h05;
            12'h1B10:q <= 8'h0E;
            12'h1B11:q <= 8'hFF;
            12'h1B12:q <= 8'h0B;
            12'h1B13:q <= 8'h0E;
            12'h1B14:q <= 8'h12;
            12'h1B15:q <= 8'hFF;
            12'h1B16:q <= 8'h0C;
            12'h1B17:q <= 8'h0D;
            12'h1B18:q <= 8'h0B;
            12'h1B19:q <= 8'hFF;
            12'h1B1A:q <= 8'h0D;
            12'h1B1B:q <= 8'h07;
            12'h1B1C:q <= 8'h0F;
            12'h1B1D:q <= 8'hFF;
            12'h1B1E:q <= 8'h0E;
            12'h1B1F:q <= 8'h03;
            12'h1B20:q <= 8'h05;
            12'h1B21:q <= 8'hFF;
            12'h1B22:q <= 8'h0F;
            12'h1B23:q <= 8'h01;
            12'h1B24:q <= 8'h03;
            12'h1B25:q <= 8'hFF;
            12'h1B26:q <= 8'h10;
            12'h1B27:q <= 8'h09;
            12'h1B28:q <= 8'h09;
            12'h1B29:q <= 8'hFF;
            12'h1B2A:q <= 8'h11;
            12'h1B2B:q <= 8'h06;
            12'h1B2C:q <= 8'h10;
            12'h1B2D:q <= 8'hFF;
            12'h1B2E:q <= 8'h12;
            12'h1B2F:q <= 8'h0C;
            12'h1B30:q <= 8'h04;
            12'h1B31:q <= 8'hFF;
            12'h1B32:q <= 8'h13;
            12'h1B33:q <= 8'h04;
            12'h1B34:q <= 8'h07;
            12'h1B35:q <= 8'hFF;
            12'h1B36:q <= 8'h00;
            12'h1B37:q <= 8'h12;
            12'h1B38:q <= 8'h0B;
            12'h1B39:q <= 8'hFF;
            12'h1B3A:q <= 8'h01;
            12'h1B3B:q <= 8'h11;
            12'h1B3C:q <= 8'h00;
            12'h1B3D:q <= 8'hFF;
            12'h1B3E:q <= 8'h02;
            12'h1B3F:q <= 8'h0A;
            12'h1B40:q <= 8'h02;
            12'h1B41:q <= 8'hFF;
            12'h1B42:q <= 8'h03;
            12'h1B43:q <= 8'h0D;
            12'h1B44:q <= 8'h04;
            12'h1B45:q <= 8'hFF;
            12'h1B46:q <= 8'h04;
            12'h1B47:q <= 8'h0E;
            12'h1B48:q <= 8'h11;
            12'h1B49:q <= 8'hFF;
            12'h1B4A:q <= 8'h05;
            12'h1B4B:q <= 8'h0F;
            12'h1B4C:q <= 8'h0A;
            12'h1B4D:q <= 8'hFF;
            12'h1B4E:q <= 8'h06;
            12'h1B4F:q <= 8'h09;
            12'h1B50:q <= 8'h10;
            12'h1B51:q <= 8'hFF;
            12'h1B52:q <= 8'h07;
            12'h1B53:q <= 8'h05;
            12'h1B54:q <= 8'h07;
            12'h1B55:q <= 8'hFF;
            12'h1B56:q <= 8'h08;
            12'h1B57:q <= 8'h02;
            12'h1B58:q <= 8'h06;
            12'h1B59:q <= 8'hFF;
            12'h1B5A:q <= 8'h09;
            12'h1B5B:q <= 8'h10;
            12'h1B5C:q <= 8'h0E;
            12'h1B5D:q <= 8'hFF;
            12'h1B5E:q <= 8'h0A;
            12'h1B5F:q <= 8'h08;
            12'h1B60:q <= 8'h13;
            12'h1B61:q <= 8'hFF;
            12'h1B62:q <= 8'h0B;
            12'h1B63:q <= 8'h07;
            12'h1B64:q <= 8'h03;
            12'h1B65:q <= 8'hFF;
            12'h1B66:q <= 8'h0C;
            12'h1B67:q <= 8'h04;
            12'h1B68:q <= 8'h0D;
            12'h1B69:q <= 8'hFF;
            12'h1B6A:q <= 8'h0D;
            12'h1B6B:q <= 8'h0C;
            12'h1B6C:q <= 8'h08;
            12'h1B6D:q <= 8'hFF;
            12'h1B6E:q <= 8'h0E;
            12'h1B6F:q <= 8'h03;
            12'h1B70:q <= 8'h09;
            12'h1B71:q <= 8'hFF;
            12'h1B72:q <= 8'h0F;
            12'h1B73:q <= 8'h06;
            12'h1B74:q <= 8'h12;
            12'h1B75:q <= 8'hFF;
            12'h1B76:q <= 8'h10;
            12'h1B77:q <= 8'h00;
            12'h1B78:q <= 8'h01;
            12'h1B79:q <= 8'hFF;
            12'h1B7A:q <= 8'h11;
            12'h1B7B:q <= 8'h01;
            12'h1B7C:q <= 8'h05;
            12'h1B7D:q <= 8'hFF;
            12'h1B7E:q <= 8'h12;
            12'h1B7F:q <= 8'h13;
            12'h1B80:q <= 8'h0F;
            12'h1B81:q <= 8'hFF;
            12'h1B82:q <= 8'h13;
            12'h1B83:q <= 8'h0B;
            12'h1B84:q <= 8'h0C;
            12'h1B85:q <= 8'hFF;
            12'h1B86:q <= 8'h00;
            12'h1B87:q <= 8'h0E;
            12'h1B88:q <= 8'h12;
            12'h1B89:q <= 8'hFF;
            12'h1B8A:q <= 8'h01;
            12'h1B8B:q <= 8'h12;
            12'h1B8C:q <= 8'h07;
            12'h1B8D:q <= 8'hFF;
            12'h1B8E:q <= 8'h02;
            12'h1B8F:q <= 8'h0B;
            12'h1B90:q <= 8'h10;
            12'h1B91:q <= 8'hFF;
            12'h1B92:q <= 8'h03;
            12'h1B93:q <= 8'h11;
            12'h1B94:q <= 8'h06;
            12'h1B95:q <= 8'hFF;
            12'h1B96:q <= 8'h04;
            12'h1B97:q <= 8'h06;
            12'h1B98:q <= 8'h05;
            12'h1B99:q <= 8'hFF;
            12'h1B9A:q <= 8'h05;
            12'h1B9B:q <= 8'h07;
            12'h1B9C:q <= 8'h03;
            12'h1B9D:q <= 8'hFF;
            12'h1B9E:q <= 8'h06;
            12'h1B9F:q <= 8'h13;
            12'h1BA0:q <= 8'h0D;
            12'h1BA1:q <= 8'hFF;
            12'h1BA2:q <= 8'h07;
            12'h1BA3:q <= 8'h0D;
            12'h1BA4:q <= 8'h0F;
            12'h1BA5:q <= 8'hFF;
            12'h1BA6:q <= 8'h08;
            12'h1BA7:q <= 8'h02;
            12'h1BA8:q <= 8'h09;
            12'h1BA9:q <= 8'hFF;
            12'h1BAA:q <= 8'h09;
            12'h1BAB:q <= 8'h04;
            12'h1BAC:q <= 8'h02;
            12'h1BAD:q <= 8'hFF;
            12'h1BAE:q <= 8'h0A;
            12'h1BAF:q <= 8'h05;
            12'h1BB0:q <= 8'h0C;
            12'h1BB1:q <= 8'hFF;
            12'h1BB2:q <= 8'h0B;
            12'h1BB3:q <= 8'h0A;
            12'h1BB4:q <= 8'h08;
            12'h1BB5:q <= 8'hFF;
            12'h1BB6:q <= 8'h0C;
            12'h1BB7:q <= 8'h0F;
            12'h1BB8:q <= 8'h00;
            12'h1BB9:q <= 8'hFF;
            12'h1BBA:q <= 8'h0D;
            12'h1BBB:q <= 8'h00;
            12'h1BBC:q <= 8'h0E;
            12'h1BBD:q <= 8'hFF;
            12'h1BBE:q <= 8'h0E;
            12'h1BBF:q <= 8'h01;
            12'h1BC0:q <= 8'h0A;
            12'h1BC1:q <= 8'hFF;
            12'h1BC2:q <= 8'h0F;
            12'h1BC3:q <= 8'h09;
            12'h1BC4:q <= 8'h11;
            12'h1BC5:q <= 8'hFF;
            12'h1BC6:q <= 8'h10;
            12'h1BC7:q <= 8'h03;
            12'h1BC8:q <= 8'h01;
            12'h1BC9:q <= 8'hFF;
            12'h1BCA:q <= 8'h11;
            12'h1BCB:q <= 8'h0C;
            12'h1BCC:q <= 8'h0B;
            12'h1BCD:q <= 8'hFF;
            12'h1BCE:q <= 8'h12;
            12'h1BCF:q <= 8'h08;
            12'h1BD0:q <= 8'h04;
            12'h1BD1:q <= 8'hFF;
            12'h1BD2:q <= 8'h13;
            12'h1BD3:q <= 8'h10;
            12'h1BD4:q <= 8'h13;
            12'h1BD5:q <= 8'hFF;
            12'h1BD6:q <= 8'h00;
            12'h1BD7:q <= 8'h03;
            12'h1BD8:q <= 8'h02;
            12'h1BD9:q <= 8'h00;
            12'h1BDA:q <= 8'hFF;
            12'h1BDB:q <= 8'h01;
            12'h1BDC:q <= 8'h00;
            12'h1BDD:q <= 8'h03;
            12'h1BDE:q <= 8'h02;
            12'h1BDF:q <= 8'hFF;
            12'h1BE0:q <= 8'h02;
            12'h1BE1:q <= 8'h01;
            12'h1BE2:q <= 8'h04;
            12'h1BE3:q <= 8'h04;
            12'h1BE4:q <= 8'hFF;
            12'h1BE5:q <= 8'h03;
            12'h1BE6:q <= 8'h04;
            12'h1BE7:q <= 8'h01;
            12'h1BE8:q <= 8'h01;
            12'h1BE9:q <= 8'hFF;
            12'h1BEA:q <= 8'h04;
            12'h1BEB:q <= 8'h02;
            12'h1BEC:q <= 8'h00;
            12'h1BED:q <= 8'h03;
            12'h1BEE:q <= 8'hFF;
            12'h1BEF:q <= 8'h00;
            12'h1BF0:q <= 8'h01;
            12'h1BF1:q <= 8'h03;
            12'h1BF2:q <= 8'hFF;
            12'h1BF3:q <= 8'h01;
            12'h1BF4:q <= 8'h02;
            12'h1BF5:q <= 8'h04;
            12'h1BF6:q <= 8'hFF;
            12'h1BF7:q <= 8'h02;
            12'h1BF8:q <= 8'h03;
            12'h1BF9:q <= 8'h01;
            12'h1BFA:q <= 8'hFF;
            12'h1BFB:q <= 8'h03;
            12'h1BFC:q <= 8'h00;
            12'h1BFD:q <= 8'h00;
            12'h1BFE:q <= 8'hFF;
            12'h1BFF:q <= 8'h04;
            12'h1C00:q <= 8'h04;
            12'h1C01:q <= 8'h02;
            12'h1C02:q <= 8'hFF;
            12'h1C03:q <= 8'h00;
            12'h1C04:q <= 8'h02;
            12'h1C05:q <= 8'h03;
            12'h1C06:q <= 8'hFF;
            12'h1C07:q <= 8'h01;
            12'h1C08:q <= 8'h03;
            12'h1C09:q <= 8'h04;
            12'h1C0A:q <= 8'hFF;
            12'h1C0B:q <= 8'h02;
            12'h1C0C:q <= 8'h04;
            12'h1C0D:q <= 8'h01;
            12'h1C0E:q <= 8'hFF;
            12'h1C0F:q <= 8'h03;
            12'h1C10:q <= 8'h00;
            12'h1C11:q <= 8'h00;
            12'h1C12:q <= 8'hFF;
            12'h1C13:q <= 8'h04;
            12'h1C14:q <= 8'h01;
            12'h1C15:q <= 8'h02;
            12'h1C16:q <= 8'hFF;
            12'h1C17:q <= 8'h00;
            12'h1C18:q <= 8'h01;
            12'h1C19:q <= 8'h01;
            12'h1C1A:q <= 8'hFF;
            12'h1C1B:q <= 8'h01;
            12'h1C1C:q <= 8'h00;
            12'h1C1D:q <= 8'h02;
            12'h1C1E:q <= 8'hFF;
            12'h1C1F:q <= 8'h02;
            12'h1C20:q <= 8'h02;
            12'h1C21:q <= 8'h03;
            12'h1C22:q <= 8'hFF;
            12'h1C23:q <= 8'h03;
            12'h1C24:q <= 8'h03;
            12'h1C25:q <= 8'h04;
            12'h1C26:q <= 8'hFF;
            12'h1C27:q <= 8'h04;
            12'h1C28:q <= 8'h04;
            12'h1C29:q <= 8'h00;
            12'h1C2A:q <= 8'hFF;
            12'h1C2B:q <= 8'h00;
            12'h1C2C:q <= 8'h04;
            12'h1C2D:q <= 8'h00;
            12'h1C2E:q <= 8'hFF;
            12'h1C2F:q <= 8'h01;
            12'h1C30:q <= 8'h02;
            12'h1C31:q <= 8'h01;
            12'h1C32:q <= 8'hFF;
            12'h1C33:q <= 8'h02;
            12'h1C34:q <= 8'h03;
            12'h1C35:q <= 8'h02;
            12'h1C36:q <= 8'hFF;
            12'h1C37:q <= 8'h03;
            12'h1C38:q <= 8'h00;
            12'h1C39:q <= 8'h03;
            12'h1C3A:q <= 8'hFF;
            12'h1C3B:q <= 8'h04;
            12'h1C3C:q <= 8'h01;
            12'h1C3D:q <= 8'h04;
            12'h1C3E:q <= 8'hFF;
            12'h1C3F:q <= 8'h00;
            12'h1C40:q <= 8'h03;
            12'h1C41:q <= 8'h02;
            12'h1C42:q <= 8'hFF;
            12'h1C43:q <= 8'h01;
            12'h1C44:q <= 8'h00;
            12'h1C45:q <= 8'h03;
            12'h1C46:q <= 8'hFF;
            12'h1C47:q <= 8'h02;
            12'h1C48:q <= 8'h01;
            12'h1C49:q <= 8'h04;
            12'h1C4A:q <= 8'hFF;
            12'h1C4B:q <= 8'h03;
            12'h1C4C:q <= 8'h04;
            12'h1C4D:q <= 8'h00;
            12'h1C4E:q <= 8'hFF;
            12'h1C4F:q <= 8'h04;
            12'h1C50:q <= 8'h02;
            12'h1C51:q <= 8'h01;
            12'h1C52:q <= 8'hFF;
            12'h1C53:q <= 8'h00;
            12'h1C54:q <= 8'h03;
            12'h1C55:q <= 8'h00;
            12'h1C56:q <= 8'hFF;
            12'h1C57:q <= 8'h01;
            12'h1C58:q <= 8'h01;
            12'h1C59:q <= 8'h04;
            12'h1C5A:q <= 8'hFF;
            12'h1C5B:q <= 8'h02;
            12'h1C5C:q <= 8'h04;
            12'h1C5D:q <= 8'h03;
            12'h1C5E:q <= 8'hFF;
            12'h1C5F:q <= 8'h03;
            12'h1C60:q <= 8'h02;
            12'h1C61:q <= 8'h02;
            12'h1C62:q <= 8'hFF;
            12'h1C63:q <= 8'h04;
            12'h1C64:q <= 8'h00;
            12'h1C65:q <= 8'h01;
            12'h1C66:q <= 8'hFF;
            12'h1C67:q <= 8'h00;
            12'h1C68:q <= 8'h01;
            12'h1C69:q <= 8'h00;
            12'h1C6A:q <= 8'hFF;
            12'h1C6B:q <= 8'h01;
            12'h1C6C:q <= 8'h02;
            12'h1C6D:q <= 8'h03;
            12'h1C6E:q <= 8'hFF;
            12'h1C6F:q <= 8'h02;
            12'h1C70:q <= 8'h03;
            12'h1C71:q <= 8'h04;
            12'h1C72:q <= 8'hFF;
            12'h1C73:q <= 8'h03;
            12'h1C74:q <= 8'h00;
            12'h1C75:q <= 8'h01;
            12'h1C76:q <= 8'hFF;
            12'h1C77:q <= 8'h04;
            12'h1C78:q <= 8'h04;
            12'h1C79:q <= 8'h02;
            12'h1C7A:q <= 8'hFF;
            12'h1C7B:q <= 8'h00;
            12'h1C7C:q <= 8'h0D;
            12'h1C7D:q <= 8'h07;
            12'h1C7E:q <= 8'h02;
            12'h1C7F:q <= 8'hFF;
            12'h1C80:q <= 8'h01;
            12'h1C81:q <= 8'h00;
            12'h1C82:q <= 8'h0B;
            12'h1C83:q <= 8'h07;
            12'h1C84:q <= 8'hFF;
            12'h1C85:q <= 8'h02;
            12'h1C86:q <= 8'h0F;
            12'h1C87:q <= 8'h06;
            12'h1C88:q <= 8'h09;
            12'h1C89:q <= 8'hFF;
            12'h1C8A:q <= 8'h03;
            12'h1C8B:q <= 8'h01;
            12'h1C8C:q <= 8'h0E;
            12'h1C8D:q <= 8'h11;
            12'h1C8E:q <= 8'hFF;
            12'h1C8F:q <= 8'h04;
            12'h1C90:q <= 8'h0B;
            12'h1C91:q <= 8'h10;
            12'h1C92:q <= 8'h04;
            12'h1C93:q <= 8'hFF;
            12'h1C94:q <= 8'h05;
            12'h1C95:q <= 8'h06;
            12'h1C96:q <= 8'h04;
            12'h1C97:q <= 8'h03;
            12'h1C98:q <= 8'hFF;
            12'h1C99:q <= 8'h06;
            12'h1C9A:q <= 8'h0C;
            12'h1C9B:q <= 8'h08;
            12'h1C9C:q <= 8'h0E;
            12'h1C9D:q <= 8'hFF;
            12'h1C9E:q <= 8'h07;
            12'h1C9F:q <= 8'h07;
            12'h1CA0:q <= 8'h0C;
            12'h1CA1:q <= 8'h01;
            12'h1CA2:q <= 8'hFF;
            12'h1CA3:q <= 8'h08;
            12'h1CA4:q <= 8'h05;
            12'h1CA5:q <= 8'h02;
            12'h1CA6:q <= 8'h06;
            12'h1CA7:q <= 8'hFF;
            12'h1CA8:q <= 8'h09;
            12'h1CA9:q <= 8'h10;
            12'h1CAA:q <= 8'h09;
            12'h1CAB:q <= 8'h0C;
            12'h1CAC:q <= 8'hFF;
            12'h1CAD:q <= 8'h0A;
            12'h1CAE:q <= 8'h0E;
            12'h1CAF:q <= 8'h11;
            12'h1CB0:q <= 8'h0A;
            12'h1CB1:q <= 8'hFF;
            12'h1CB2:q <= 8'h0B;
            12'h1CB3:q <= 8'h08;
            12'h1CB4:q <= 8'h05;
            12'h1CB5:q <= 8'h00;
            12'h1CB6:q <= 8'hFF;
            12'h1CB7:q <= 8'h0C;
            12'h1CB8:q <= 8'h03;
            12'h1CB9:q <= 8'h01;
            12'h1CBA:q <= 8'h0B;
            12'h1CBB:q <= 8'hFF;
            12'h1CBC:q <= 8'h0D;
            12'h1CBD:q <= 8'h11;
            12'h1CBE:q <= 8'h00;
            12'h1CBF:q <= 8'h0F;
            12'h1CC0:q <= 8'hFF;
            12'h1CC1:q <= 8'h0E;
            12'h1CC2:q <= 8'h04;
            12'h1CC3:q <= 8'h0A;
            12'h1CC4:q <= 8'h10;
            12'h1CC5:q <= 8'hFF;
            12'h1CC6:q <= 8'h0F;
            12'h1CC7:q <= 8'h09;
            12'h1CC8:q <= 8'h0D;
            12'h1CC9:q <= 8'h0D;
            12'h1CCA:q <= 8'hFF;
            12'h1CCB:q <= 8'h10;
            12'h1CCC:q <= 8'h02;
            12'h1CCD:q <= 8'h03;
            12'h1CCE:q <= 8'h05;
            12'h1CCF:q <= 8'hFF;
            12'h1CD0:q <= 8'h11;
            12'h1CD1:q <= 8'h0A;
            12'h1CD2:q <= 8'h0F;
            12'h1CD3:q <= 8'h08;
            12'h1CD4:q <= 8'hFF;
            12'h1CD5:q <= 8'h00;
            12'h1CD6:q <= 8'h10;
            12'h1CD7:q <= 8'h05;
            12'h1CD8:q <= 8'hFF;
            12'h1CD9:q <= 8'h01;
            12'h1CDA:q <= 8'h06;
            12'h1CDB:q <= 8'h0E;
            12'h1CDC:q <= 8'hFF;
            12'h1CDD:q <= 8'h02;
            12'h1CDE:q <= 8'h03;
            12'h1CDF:q <= 8'h0D;
            12'h1CE0:q <= 8'hFF;
            12'h1CE1:q <= 8'h03;
            12'h1CE2:q <= 8'h0E;
            12'h1CE3:q <= 8'h06;
            12'h1CE4:q <= 8'hFF;
            12'h1CE5:q <= 8'h04;
            12'h1CE6:q <= 8'h04;
            12'h1CE7:q <= 8'h0F;
            12'h1CE8:q <= 8'hFF;
            12'h1CE9:q <= 8'h05;
            12'h1CEA:q <= 8'h09;
            12'h1CEB:q <= 8'h03;
            12'h1CEC:q <= 8'hFF;
            12'h1CED:q <= 8'h06;
            12'h1CEE:q <= 8'h07;
            12'h1CEF:q <= 8'h04;
            12'h1CF0:q <= 8'hFF;
            12'h1CF1:q <= 8'h07;
            12'h1CF2:q <= 8'h11;
            12'h1CF3:q <= 8'h11;
            12'h1CF4:q <= 8'hFF;
            12'h1CF5:q <= 8'h08;
            12'h1CF6:q <= 8'h00;
            12'h1CF7:q <= 8'h08;
            12'h1CF8:q <= 8'hFF;
            12'h1CF9:q <= 8'h09;
            12'h1CFA:q <= 8'h02;
            12'h1CFB:q <= 8'h09;
            12'h1CFC:q <= 8'hFF;
            12'h1CFD:q <= 8'h0A;
            12'h1CFE:q <= 8'h0F;
            12'h1CFF:q <= 8'h07;
            12'h1D00:q <= 8'hFF;
            12'h1D01:q <= 8'h0B;
            12'h1D02:q <= 8'h0D;
            12'h1D03:q <= 8'h0B;
            12'h1D04:q <= 8'hFF;
            12'h1D05:q <= 8'h0C;
            12'h1D06:q <= 8'h08;
            12'h1D07:q <= 8'h01;
            12'h1D08:q <= 8'hFF;
            12'h1D09:q <= 8'h0D;
            12'h1D0A:q <= 8'h01;
            12'h1D0B:q <= 8'h0C;
            12'h1D0C:q <= 8'hFF;
            12'h1D0D:q <= 8'h0E;
            12'h1D0E:q <= 8'h05;
            12'h1D0F:q <= 8'h0A;
            12'h1D10:q <= 8'hFF;
            12'h1D11:q <= 8'h0F;
            12'h1D12:q <= 8'h0A;
            12'h1D13:q <= 8'h10;
            12'h1D14:q <= 8'hFF;
            12'h1D15:q <= 8'h10;
            12'h1D16:q <= 8'h0B;
            12'h1D17:q <= 8'h02;
            12'h1D18:q <= 8'hFF;
            12'h1D19:q <= 8'h11;
            12'h1D1A:q <= 8'h0C;
            12'h1D1B:q <= 8'h00;
            12'h1D1C:q <= 8'hFF;
            12'h1D1D:q <= 8'h00;
            12'h1D1E:q <= 8'h07;
            12'h1D1F:q <= 8'h02;
            12'h1D20:q <= 8'hFF;
            12'h1D21:q <= 8'h01;
            12'h1D22:q <= 8'h10;
            12'h1D23:q <= 8'h00;
            12'h1D24:q <= 8'hFF;
            12'h1D25:q <= 8'h02;
            12'h1D26:q <= 8'h0A;
            12'h1D27:q <= 8'h0B;
            12'h1D28:q <= 8'hFF;
            12'h1D29:q <= 8'h03;
            12'h1D2A:q <= 8'h03;
            12'h1D2B:q <= 8'h11;
            12'h1D2C:q <= 8'hFF;
            12'h1D2D:q <= 8'h04;
            12'h1D2E:q <= 8'h02;
            12'h1D2F:q <= 8'h06;
            12'h1D30:q <= 8'hFF;
            12'h1D31:q <= 8'h05;
            12'h1D32:q <= 8'h0E;
            12'h1D33:q <= 8'h07;
            12'h1D34:q <= 8'hFF;
            12'h1D35:q <= 8'h06;
            12'h1D36:q <= 8'h0C;
            12'h1D37:q <= 8'h09;
            12'h1D38:q <= 8'hFF;
            12'h1D39:q <= 8'h07;
            12'h1D3A:q <= 8'h09;
            12'h1D3B:q <= 8'h0D;
            12'h1D3C:q <= 8'hFF;
            12'h1D3D:q <= 8'h08;
            12'h1D3E:q <= 8'h01;
            12'h1D3F:q <= 8'h01;
            12'h1D40:q <= 8'hFF;
            12'h1D41:q <= 8'h09;
            12'h1D42:q <= 8'h0D;
            12'h1D43:q <= 8'h04;
            12'h1D44:q <= 8'hFF;
            12'h1D45:q <= 8'h0A;
            12'h1D46:q <= 8'h05;
            12'h1D47:q <= 8'h05;
            12'h1D48:q <= 8'hFF;
            12'h1D49:q <= 8'h0B;
            12'h1D4A:q <= 8'h08;
            12'h1D4B:q <= 8'h08;
            12'h1D4C:q <= 8'hFF;
            12'h1D4D:q <= 8'h0C;
            12'h1D4E:q <= 8'h0B;
            12'h1D4F:q <= 8'h0E;
            12'h1D50:q <= 8'hFF;
            12'h1D51:q <= 8'h0D;
            12'h1D52:q <= 8'h0F;
            12'h1D53:q <= 8'h0F;
            12'h1D54:q <= 8'hFF;
            12'h1D55:q <= 8'h0E;
            12'h1D56:q <= 8'h11;
            12'h1D57:q <= 8'h0C;
            12'h1D58:q <= 8'hFF;
            12'h1D59:q <= 8'h0F;
            12'h1D5A:q <= 8'h04;
            12'h1D5B:q <= 8'h0A;
            12'h1D5C:q <= 8'hFF;
            12'h1D5D:q <= 8'h10;
            12'h1D5E:q <= 8'h06;
            12'h1D5F:q <= 8'h03;
            12'h1D60:q <= 8'hFF;
            12'h1D61:q <= 8'h11;
            12'h1D62:q <= 8'h00;
            12'h1D63:q <= 8'h10;
            12'h1D64:q <= 8'hFF;
            12'h1D65:q <= 8'h00;
            12'h1D66:q <= 8'h0A;
            12'h1D67:q <= 8'h11;
            12'h1D68:q <= 8'hFF;
            12'h1D69:q <= 8'h01;
            12'h1D6A:q <= 8'h08;
            12'h1D6B:q <= 8'h0B;
            12'h1D6C:q <= 8'hFF;
            12'h1D6D:q <= 8'h02;
            12'h1D6E:q <= 8'h07;
            12'h1D6F:q <= 8'h01;
            12'h1D70:q <= 8'hFF;
            12'h1D71:q <= 8'h03;
            12'h1D72:q <= 8'h0D;
            12'h1D73:q <= 8'h00;
            12'h1D74:q <= 8'hFF;
            12'h1D75:q <= 8'h04;
            12'h1D76:q <= 8'h02;
            12'h1D77:q <= 8'h07;
            12'h1D78:q <= 8'hFF;
            12'h1D79:q <= 8'h05;
            12'h1D7A:q <= 8'h05;
            12'h1D7B:q <= 8'h10;
            12'h1D7C:q <= 8'hFF;
            12'h1D7D:q <= 8'h06;
            12'h1D7E:q <= 8'h09;
            12'h1D7F:q <= 8'h06;
            12'h1D80:q <= 8'hFF;
            12'h1D81:q <= 8'h07;
            12'h1D82:q <= 8'h04;
            12'h1D83:q <= 8'h05;
            12'h1D84:q <= 8'hFF;
            12'h1D85:q <= 8'h08;
            12'h1D86:q <= 8'h01;
            12'h1D87:q <= 8'h02;
            12'h1D88:q <= 8'hFF;
            12'h1D89:q <= 8'h09;
            12'h1D8A:q <= 8'h0F;
            12'h1D8B:q <= 8'h08;
            12'h1D8C:q <= 8'hFF;
            12'h1D8D:q <= 8'h0A;
            12'h1D8E:q <= 8'h00;
            12'h1D8F:q <= 8'h0C;
            12'h1D90:q <= 8'hFF;
            12'h1D91:q <= 8'h0B;
            12'h1D92:q <= 8'h10;
            12'h1D93:q <= 8'h0E;
            12'h1D94:q <= 8'hFF;
            12'h1D95:q <= 8'h0C;
            12'h1D96:q <= 8'h0C;
            12'h1D97:q <= 8'h0F;
            12'h1D98:q <= 8'hFF;
            12'h1D99:q <= 8'h0D;
            12'h1D9A:q <= 8'h0B;
            12'h1D9B:q <= 8'h0A;
            12'h1D9C:q <= 8'hFF;
            12'h1D9D:q <= 8'h0E;
            12'h1D9E:q <= 8'h06;
            12'h1D9F:q <= 8'h04;
            12'h1DA0:q <= 8'hFF;
            12'h1DA1:q <= 8'h0F;
            12'h1DA2:q <= 8'h03;
            12'h1DA3:q <= 8'h0D;
            12'h1DA4:q <= 8'hFF;
            12'h1DA5:q <= 8'h10;
            12'h1DA6:q <= 8'h0E;
            12'h1DA7:q <= 8'h09;
            12'h1DA8:q <= 8'hFF;
            12'h1DA9:q <= 8'h11;
            12'h1DAA:q <= 8'h11;
            12'h1DAB:q <= 8'h03;
            12'h1DAC:q <= 8'hFF;
            12'h1DAD:q <= 8'h00;
            12'h1DAE:q <= 8'h09;
            12'h1DAF:q <= 8'h0B;
            12'h1DB0:q <= 8'hFF;
            12'h1DB1:q <= 8'h01;
            12'h1DB2:q <= 8'h0B;
            12'h1DB3:q <= 8'h0A;
            12'h1DB4:q <= 8'hFF;
            12'h1DB5:q <= 8'h02;
            12'h1DB6:q <= 8'h05;
            12'h1DB7:q <= 8'h05;
            12'h1DB8:q <= 8'hFF;
            12'h1DB9:q <= 8'h03;
            12'h1DBA:q <= 8'h0E;
            12'h1DBB:q <= 8'h01;
            12'h1DBC:q <= 8'hFF;
            12'h1DBD:q <= 8'h04;
            12'h1DBE:q <= 8'h0C;
            12'h1DBF:q <= 8'h10;
            12'h1DC0:q <= 8'hFF;
            12'h1DC1:q <= 8'h05;
            12'h1DC2:q <= 8'h10;
            12'h1DC3:q <= 8'h04;
            12'h1DC4:q <= 8'hFF;
            12'h1DC5:q <= 8'h06;
            12'h1DC6:q <= 8'h06;
            12'h1DC7:q <= 8'h03;
            12'h1DC8:q <= 8'hFF;
            12'h1DC9:q <= 8'h07;
            12'h1DCA:q <= 8'h03;
            12'h1DCB:q <= 8'h02;
            12'h1DCC:q <= 8'hFF;
            12'h1DCD:q <= 8'h08;
            12'h1DCE:q <= 8'h04;
            12'h1DCF:q <= 8'h09;
            12'h1DD0:q <= 8'hFF;
            12'h1DD1:q <= 8'h09;
            12'h1DD2:q <= 8'h07;
            12'h1DD3:q <= 8'h0E;
            12'h1DD4:q <= 8'hFF;
            12'h1DD5:q <= 8'h0A;
            12'h1DD6:q <= 8'h02;
            12'h1DD7:q <= 8'h0D;
            12'h1DD8:q <= 8'hFF;
            12'h1DD9:q <= 8'h0B;
            12'h1DDA:q <= 8'h0F;
            12'h1DDB:q <= 8'h0C;
            12'h1DDC:q <= 8'hFF;
            12'h1DDD:q <= 8'h0C;
            12'h1DDE:q <= 8'h00;
            12'h1DDF:q <= 8'h07;
            12'h1DE0:q <= 8'hFF;
            12'h1DE1:q <= 8'h0D;
            12'h1DE2:q <= 8'h0D;
            12'h1DE3:q <= 8'h0F;
            12'h1DE4:q <= 8'hFF;
            12'h1DE5:q <= 8'h0E;
            12'h1DE6:q <= 8'h11;
            12'h1DE7:q <= 8'h00;
            12'h1DE8:q <= 8'hFF;
            12'h1DE9:q <= 8'h0F;
            12'h1DEA:q <= 8'h01;
            12'h1DEB:q <= 8'h06;
            12'h1DEC:q <= 8'hFF;
            12'h1DED:q <= 8'h10;
            12'h1DEE:q <= 8'h08;
            12'h1DEF:q <= 8'h08;
            12'h1DF0:q <= 8'hFF;
            12'h1DF1:q <= 8'h11;
            12'h1DF2:q <= 8'h0A;
            12'h1DF3:q <= 8'h11;
            12'h1DF4:q <= 8'hFF;
            12'h1DF5:q <= 8'h00;
            12'h1DF6:q <= 8'h04;
            12'h1DF7:q <= 8'h04;
            12'h1DF8:q <= 8'hFF;
            12'h1DF9:q <= 8'h01;
            12'h1DFA:q <= 8'h07;
            12'h1DFB:q <= 8'h00;
            12'h1DFC:q <= 8'hFF;
            12'h1DFD:q <= 8'h02;
            12'h1DFE:q <= 8'h05;
            12'h1DFF:q <= 8'h07;
            12'h1E00:q <= 8'hFF;
            12'h1E01:q <= 8'h03;
            12'h1E02:q <= 8'h06;
            12'h1E03:q <= 8'h0A;
            12'h1E04:q <= 8'hFF;
            12'h1E05:q <= 8'h04;
            12'h1E06:q <= 8'h01;
            12'h1E07:q <= 8'h11;
            12'h1E08:q <= 8'hFF;
            12'h1E09:q <= 8'h05;
            12'h1E0A:q <= 8'h0E;
            12'h1E0B:q <= 8'h06;
            12'h1E0C:q <= 8'hFF;
            12'h1E0D:q <= 8'h06;
            12'h1E0E:q <= 8'h11;
            12'h1E0F:q <= 8'h0C;
            12'h1E10:q <= 8'hFF;
            12'h1E11:q <= 8'h07;
            12'h1E12:q <= 8'h00;
            12'h1E13:q <= 8'h09;
            12'h1E14:q <= 8'hFF;
            12'h1E15:q <= 8'h08;
            12'h1E16:q <= 8'h10;
            12'h1E17:q <= 8'h02;
            12'h1E18:q <= 8'hFF;
            12'h1E19:q <= 8'h09;
            12'h1E1A:q <= 8'h0F;
            12'h1E1B:q <= 8'h0E;
            12'h1E1C:q <= 8'hFF;
            12'h1E1D:q <= 8'h0A;
            12'h1E1E:q <= 8'h02;
            12'h1E1F:q <= 8'h01;
            12'h1E20:q <= 8'hFF;
            12'h1E21:q <= 8'h0B;
            12'h1E22:q <= 8'h0B;
            12'h1E23:q <= 8'h0D;
            12'h1E24:q <= 8'hFF;
            12'h1E25:q <= 8'h0C;
            12'h1E26:q <= 8'h08;
            12'h1E27:q <= 8'h0B;
            12'h1E28:q <= 8'hFF;
            12'h1E29:q <= 8'h0D;
            12'h1E2A:q <= 8'h0D;
            12'h1E2B:q <= 8'h10;
            12'h1E2C:q <= 8'hFF;
            12'h1E2D:q <= 8'h0E;
            12'h1E2E:q <= 8'h0A;
            12'h1E2F:q <= 8'h0F;
            12'h1E30:q <= 8'hFF;
            12'h1E31:q <= 8'h0F;
            12'h1E32:q <= 8'h03;
            12'h1E33:q <= 8'h05;
            12'h1E34:q <= 8'hFF;
            12'h1E35:q <= 8'h10;
            12'h1E36:q <= 8'h09;
            12'h1E37:q <= 8'h03;
            12'h1E38:q <= 8'hFF;
            12'h1E39:q <= 8'h11;
            12'h1E3A:q <= 8'h0C;
            12'h1E3B:q <= 8'h08;
            12'h1E3C:q <= 8'hFF;
            12'h1E3D:q <= 8'h00;
            12'h1E3E:q <= 8'h03;
            12'h1E3F:q <= 8'h0A;
            12'h1E40:q <= 8'hFF;
            12'h1E41:q <= 8'h01;
            12'h1E42:q <= 8'h02;
            12'h1E43:q <= 8'h08;
            12'h1E44:q <= 8'hFF;
            12'h1E45:q <= 8'h02;
            12'h1E46:q <= 8'h0C;
            12'h1E47:q <= 8'h03;
            12'h1E48:q <= 8'hFF;
            12'h1E49:q <= 8'h03;
            12'h1E4A:q <= 8'h10;
            12'h1E4B:q <= 8'h0B;
            12'h1E4C:q <= 8'hFF;
            12'h1E4D:q <= 8'h04;
            12'h1E4E:q <= 8'h0F;
            12'h1E4F:q <= 8'h00;
            12'h1E50:q <= 8'hFF;
            12'h1E51:q <= 8'h05;
            12'h1E52:q <= 8'h0E;
            12'h1E53:q <= 8'h06;
            12'h1E54:q <= 8'hFF;
            12'h1E55:q <= 8'h06;
            12'h1E56:q <= 8'h0A;
            12'h1E57:q <= 8'h04;
            12'h1E58:q <= 8'hFF;
            12'h1E59:q <= 8'h07;
            12'h1E5A:q <= 8'h04;
            12'h1E5B:q <= 8'h0F;
            12'h1E5C:q <= 8'hFF;
            12'h1E5D:q <= 8'h08;
            12'h1E5E:q <= 8'h07;
            12'h1E5F:q <= 8'h07;
            12'h1E60:q <= 8'hFF;
            12'h1E61:q <= 8'h09;
            12'h1E62:q <= 8'h11;
            12'h1E63:q <= 8'h0D;
            12'h1E64:q <= 8'hFF;
            12'h1E65:q <= 8'h0A;
            12'h1E66:q <= 8'h08;
            12'h1E67:q <= 8'h01;
            12'h1E68:q <= 8'hFF;
            12'h1E69:q <= 8'h0B;
            12'h1E6A:q <= 8'h01;
            12'h1E6B:q <= 8'h0C;
            12'h1E6C:q <= 8'hFF;
            12'h1E6D:q <= 8'h0C;
            12'h1E6E:q <= 8'h0B;
            12'h1E6F:q <= 8'h09;
            12'h1E70:q <= 8'hFF;
            12'h1E71:q <= 8'h0D;
            12'h1E72:q <= 8'h06;
            12'h1E73:q <= 8'h05;
            12'h1E74:q <= 8'hFF;
            12'h1E75:q <= 8'h0E;
            12'h1E76:q <= 8'h05;
            12'h1E77:q <= 8'h0E;
            12'h1E78:q <= 8'hFF;
            12'h1E79:q <= 8'h0F;
            12'h1E7A:q <= 8'h09;
            12'h1E7B:q <= 8'h11;
            12'h1E7C:q <= 8'hFF;
            12'h1E7D:q <= 8'h10;
            12'h1E7E:q <= 8'h00;
            12'h1E7F:q <= 8'h02;
            12'h1E80:q <= 8'hFF;
            12'h1E81:q <= 8'h11;
            12'h1E82:q <= 8'h0D;
            12'h1E83:q <= 8'h10;
            12'h1E84:q <= 8'hFF;
            12'h1E85:q <= 8'h00;
            12'h1E86:q <= 8'h04;
            12'h1E87:q <= 8'h00;
            12'h1E88:q <= 8'hFF;
            12'h1E89:q <= 8'h01;
            12'h1E8A:q <= 8'h0E;
            12'h1E8B:q <= 8'h10;
            12'h1E8C:q <= 8'hFF;
            12'h1E8D:q <= 8'h02;
            12'h1E8E:q <= 8'h0F;
            12'h1E8F:q <= 8'h09;
            12'h1E90:q <= 8'hFF;
            12'h1E91:q <= 8'h03;
            12'h1E92:q <= 8'h0C;
            12'h1E93:q <= 8'h0F;
            12'h1E94:q <= 8'hFF;
            12'h1E95:q <= 8'h04;
            12'h1E96:q <= 8'h0B;
            12'h1E97:q <= 8'h0C;
            12'h1E98:q <= 8'hFF;
            12'h1E99:q <= 8'h05;
            12'h1E9A:q <= 8'h00;
            12'h1E9B:q <= 8'h08;
            12'h1E9C:q <= 8'hFF;
            12'h1E9D:q <= 8'h06;
            12'h1E9E:q <= 8'h05;
            12'h1E9F:q <= 8'h0A;
            12'h1EA0:q <= 8'hFF;
            12'h1EA1:q <= 8'h07;
            12'h1EA2:q <= 8'h11;
            12'h1EA3:q <= 8'h05;
            12'h1EA4:q <= 8'hFF;
            12'h1EA5:q <= 8'h08;
            12'h1EA6:q <= 8'h07;
            12'h1EA7:q <= 8'h04;
            12'h1EA8:q <= 8'hFF;
            12'h1EA9:q <= 8'h09;
            12'h1EAA:q <= 8'h06;
            12'h1EAB:q <= 8'h03;
            12'h1EAC:q <= 8'hFF;
            12'h1EAD:q <= 8'h0A;
            12'h1EAE:q <= 8'h0D;
            12'h1EAF:q <= 8'h07;
            12'h1EB0:q <= 8'hFF;
            12'h1EB1:q <= 8'h0B;
            12'h1EB2:q <= 8'h02;
            12'h1EB3:q <= 8'h0B;
            12'h1EB4:q <= 8'hFF;
            12'h1EB5:q <= 8'h0C;
            12'h1EB6:q <= 8'h03;
            12'h1EB7:q <= 8'h0D;
            12'h1EB8:q <= 8'hFF;
            12'h1EB9:q <= 8'h0D;
            12'h1EBA:q <= 8'h0A;
            12'h1EBB:q <= 8'h06;
            12'h1EBC:q <= 8'hFF;
            12'h1EBD:q <= 8'h0E;
            12'h1EBE:q <= 8'h09;
            12'h1EBF:q <= 8'h01;
            12'h1EC0:q <= 8'hFF;
            12'h1EC1:q <= 8'h0F;
            12'h1EC2:q <= 8'h08;
            12'h1EC3:q <= 8'h11;
            12'h1EC4:q <= 8'hFF;
            12'h1EC5:q <= 8'h10;
            12'h1EC6:q <= 8'h10;
            12'h1EC7:q <= 8'h0E;
            12'h1EC8:q <= 8'hFF;
            12'h1EC9:q <= 8'h11;
            12'h1ECA:q <= 8'h01;
            12'h1ECB:q <= 8'h02;
            12'h1ECC:q <= 8'hFF;
            12'h1ECD:q <= 8'h00;
            12'h1ECE:q <= 8'h01;
            12'h1ECF:q <= 8'h0C;
            12'h1ED0:q <= 8'hFF;
            12'h1ED1:q <= 8'h01;
            12'h1ED2:q <= 8'h09;
            12'h1ED3:q <= 8'h0D;
            12'h1ED4:q <= 8'hFF;
            12'h1ED5:q <= 8'h02;
            12'h1ED6:q <= 8'h03;
            12'h1ED7:q <= 8'h02;
            12'h1ED8:q <= 8'hFF;
            12'h1ED9:q <= 8'h03;
            12'h1EDA:q <= 8'h0B;
            12'h1EDB:q <= 8'h0E;
            12'h1EDC:q <= 8'hFF;
            12'h1EDD:q <= 8'h04;
            12'h1EDE:q <= 8'h07;
            12'h1EDF:q <= 8'h06;
            12'h1EE0:q <= 8'hFF;
            12'h1EE1:q <= 8'h05;
            12'h1EE2:q <= 8'h05;
            12'h1EE3:q <= 8'h10;
            12'h1EE4:q <= 8'hFF;
            12'h1EE5:q <= 8'h06;
            12'h1EE6:q <= 8'h10;
            12'h1EE7:q <= 8'h08;
            12'h1EE8:q <= 8'hFF;
            12'h1EE9:q <= 8'h07;
            12'h1EEA:q <= 8'h06;
            12'h1EEB:q <= 8'h0F;
            12'h1EEC:q <= 8'hFF;
            12'h1EED:q <= 8'h08;
            12'h1EEE:q <= 8'h04;
            12'h1EEF:q <= 8'h03;
            12'h1EF0:q <= 8'hFF;
            12'h1EF1:q <= 8'h09;
            12'h1EF2:q <= 8'h0E;
            12'h1EF3:q <= 8'h00;
            12'h1EF4:q <= 8'hFF;
            12'h1EF5:q <= 8'h0A;
            12'h1EF6:q <= 8'h00;
            12'h1EF7:q <= 8'h0A;
            12'h1EF8:q <= 8'hFF;
            12'h1EF9:q <= 8'h0B;
            12'h1EFA:q <= 8'h0F;
            12'h1EFB:q <= 8'h04;
            12'h1EFC:q <= 8'hFF;
            12'h1EFD:q <= 8'h0C;
            12'h1EFE:q <= 8'h11;
            12'h1EFF:q <= 8'h07;
            12'h1F00:q <= 8'hFF;
            12'h1F01:q <= 8'h0D;
            12'h1F02:q <= 8'h0D;
            12'h1F03:q <= 8'h11;
            12'h1F04:q <= 8'hFF;
            12'h1F05:q <= 8'h0E;
            12'h1F06:q <= 8'h0C;
            12'h1F07:q <= 8'h01;
            12'h1F08:q <= 8'hFF;
            12'h1F09:q <= 8'h0F;
            12'h1F0A:q <= 8'h02;
            12'h1F0B:q <= 8'h05;
            12'h1F0C:q <= 8'hFF;
            12'h1F0D:q <= 8'h10;
            12'h1F0E:q <= 8'h0A;
            12'h1F0F:q <= 8'h09;
            12'h1F10:q <= 8'hFF;
            12'h1F11:q <= 8'h11;
            12'h1F12:q <= 8'h08;
            12'h1F13:q <= 8'h0B;
            12'h1F14:q <= 8'hFF;
            12'h1F15:q <= 8'h00;
            12'h1F16:q <= 8'h00;
            12'h1F17:q <= 8'h00;
            12'h1F18:q <= 8'h00;
            12'h1F19:q <= 8'h00;
            12'h1F1A:q <= 8'h00;
            12'h1F1B:q <= 8'h00;
            12'h1F1C:q <= 8'h00;
            12'h1F1D:q <= 8'h00;
            12'h1F1E:q <= 8'h00;
            12'h1F1F:q <= 8'h00;
            12'h1F20:q <= 8'h00;
            12'h1F21:q <= 8'h00;
            12'h1F22:q <= 8'h00;
            12'h1F23:q <= 8'h00;
            12'h1F24:q <= 8'h00;
            12'h1F25:q <= 8'h00;
            12'h1F26:q <= 8'h00;
            12'h1F27:q <= 8'h00;
            12'h1F28:q <= 8'h00;
            12'h1F29:q <= 8'h00;
            12'h1F2A:q <= 8'h00;
            12'h1F2B:q <= 8'h00;
            12'h1F2C:q <= 8'h00;
            12'h1F2D:q <= 8'h00;
            12'h1F2E:q <= 8'h00;
            12'h1F2F:q <= 8'h00;
            12'h1F30:q <= 8'h00;
            12'h1F31:q <= 8'h00;
            12'h1F32:q <= 8'h00;
            12'h1F33:q <= 8'h00;
            12'h1F34:q <= 8'h00;
            12'h1F35:q <= 8'h00;
            12'h1F36:q <= 8'h00;
            12'h1F37:q <= 8'h00;
            12'h1F38:q <= 8'h00;
            12'h1F39:q <= 8'h00;
            12'h1F3A:q <= 8'h00;
            12'h1F3B:q <= 8'h00;
            12'h1F3C:q <= 8'h00;
            12'h1F3D:q <= 8'h00;
            12'h1F3E:q <= 8'h00;
            12'h1F3F:q <= 8'h00;
            12'h1F40:q <= 8'h00;
            12'h1F41:q <= 8'h00;
            12'h1F42:q <= 8'h00;
            12'h1F43:q <= 8'h00;
            12'h1F44:q <= 8'h00;
            12'h1F45:q <= 8'h00;
            12'h1F46:q <= 8'h00;
            12'h1F47:q <= 8'h00;
            12'h1F48:q <= 8'h00;
            12'h1F49:q <= 8'h00;
            12'h1F4A:q <= 8'h00;
            12'h1F4B:q <= 8'h00;
            12'h1F4C:q <= 8'h00;
            12'h1F4D:q <= 8'h00;
            12'h1F4E:q <= 8'h00;
            12'h1F4F:q <= 8'h00;
            12'h1F50:q <= 8'h00;
            12'h1F51:q <= 8'h00;
            12'h1F52:q <= 8'h00;
            12'h1F53:q <= 8'h00;
            12'h1F54:q <= 8'h00;
            12'h1F55:q <= 8'h00;
            12'h1F56:q <= 8'h00;
            12'h1F57:q <= 8'h00;
            12'h1F58:q <= 8'h00;
            12'h1F59:q <= 8'h00;
            12'h1F5A:q <= 8'h00;
            12'h1F5B:q <= 8'h00;
            12'h1F5C:q <= 8'h00;
            12'h1F5D:q <= 8'h00;
            12'h1F5E:q <= 8'h00;
            12'h1F5F:q <= 8'h00;
            12'h1F60:q <= 8'h00;
            12'h1F61:q <= 8'h00;
            12'h1F62:q <= 8'h00;
            12'h1F63:q <= 8'h00;
            12'h1F64:q <= 8'h00;
            12'h1F65:q <= 8'h00;
            12'h1F66:q <= 8'h00;
            12'h1F67:q <= 8'h00;
            12'h1F68:q <= 8'h00;
            12'h1F69:q <= 8'h00;
            12'h1F6A:q <= 8'h00;
            12'h1F6B:q <= 8'h00;
            12'h1F6C:q <= 8'h00;
            12'h1F6D:q <= 8'h00;
            12'h1F6E:q <= 8'h00;
            12'h1F6F:q <= 8'h00;
            12'h1F70:q <= 8'h00;
            12'h1F71:q <= 8'h00;
            12'h1F72:q <= 8'h00;
            12'h1F73:q <= 8'h00;
            12'h1F74:q <= 8'h00;
            12'h1F75:q <= 8'h00;
            12'h1F76:q <= 8'h00;
            12'h1F77:q <= 8'h00;
            12'h1F78:q <= 8'h00;
            12'h1F79:q <= 8'h00;
            12'h1F7A:q <= 8'h00;
            12'h1F7B:q <= 8'h00;
            12'h1F7C:q <= 8'h00;
            12'h1F7D:q <= 8'h00;
            12'h1F7E:q <= 8'h00;
            12'h1F7F:q <= 8'h00;
            12'h1F80:q <= 8'h00;
            12'h1F81:q <= 8'h00;
            12'h1F82:q <= 8'h00;
            12'h1F83:q <= 8'h00;
            12'h1F84:q <= 8'h00;
            12'h1F85:q <= 8'h00;
            12'h1F86:q <= 8'h00;
            12'h1F87:q <= 8'h00;
            12'h1F88:q <= 8'h00;
            12'h1F89:q <= 8'h00;
            12'h1F8A:q <= 8'h00;
            12'h1F8B:q <= 8'h00;
            12'h1F8C:q <= 8'h00;
            12'h1F8D:q <= 8'h00;
            12'h1F8E:q <= 8'h00;
            12'h1F8F:q <= 8'h00;
            12'h1F90:q <= 8'h00;
            12'h1F91:q <= 8'h00;
            12'h1F92:q <= 8'h00;
            12'h1F93:q <= 8'h00;
            12'h1F94:q <= 8'h00;
            12'h1F95:q <= 8'h00;
            12'h1F96:q <= 8'h00;
            12'h1F97:q <= 8'h00;
            12'h1F98:q <= 8'h00;
            12'h1F99:q <= 8'h00;
            12'h1F9A:q <= 8'h00;
            12'h1F9B:q <= 8'h00;
            12'h1F9C:q <= 8'h00;
            12'h1F9D:q <= 8'h00;
            12'h1F9E:q <= 8'h00;
            12'h1F9F:q <= 8'h00;
            12'h1FA0:q <= 8'h00;
            12'h1FA1:q <= 8'h00;
            12'h1FA2:q <= 8'h00;
            12'h1FA3:q <= 8'h00;
            12'h1FA4:q <= 8'h00;
            12'h1FA5:q <= 8'h00;
            12'h1FA6:q <= 8'h00;
            12'h1FA7:q <= 8'h00;
            12'h1FA8:q <= 8'h00;
            12'h1FA9:q <= 8'h00;
            12'h1FAA:q <= 8'h00;
            12'h1FAB:q <= 8'h00;
            12'h1FAC:q <= 8'h00;
            12'h1FAD:q <= 8'h00;
            12'h1FAE:q <= 8'h00;
            12'h1FAF:q <= 8'h00;
            12'h1FB0:q <= 8'h00;
            12'h1FB1:q <= 8'h00;
            12'h1FB2:q <= 8'h00;
            12'h1FB3:q <= 8'h00;
            12'h1FB4:q <= 8'h00;
            12'h1FB5:q <= 8'h00;
            12'h1FB6:q <= 8'h00;
            12'h1FB7:q <= 8'h00;
            12'h1FB8:q <= 8'h00;
            12'h1FB9:q <= 8'h00;
            12'h1FBA:q <= 8'h00;
            12'h1FBB:q <= 8'h00;
            12'h1FBC:q <= 8'h00;
            12'h1FBD:q <= 8'h00;
            12'h1FBE:q <= 8'h00;
            12'h1FBF:q <= 8'h00;
            12'h1FC0:q <= 8'h00;
            12'h1FC1:q <= 8'h00;
            12'h1FC2:q <= 8'h00;
            12'h1FC3:q <= 8'h00;
            12'h1FC4:q <= 8'h00;
            12'h1FC5:q <= 8'h00;
            12'h1FC6:q <= 8'h00;
            12'h1FC7:q <= 8'h00;
            12'h1FC8:q <= 8'h00;
            12'h1FC9:q <= 8'h00;
            12'h1FCA:q <= 8'h00;
            12'h1FCB:q <= 8'h00;
            12'h1FCC:q <= 8'h00;
            12'h1FCD:q <= 8'h00;
            12'h1FCE:q <= 8'h00;
            12'h1FCF:q <= 8'h00;
            12'h1FD0:q <= 8'h00;
            12'h1FD1:q <= 8'h00;
            12'h1FD2:q <= 8'h00;
            12'h1FD3:q <= 8'h00;
            12'h1FD4:q <= 8'h00;
            12'h1FD5:q <= 8'h00;
            12'h1FD6:q <= 8'h00;
            12'h1FD7:q <= 8'h00;
            12'h1FD8:q <= 8'h00;
            12'h1FD9:q <= 8'h00;
            12'h1FDA:q <= 8'h00;
            12'h1FDB:q <= 8'h00;
            12'h1FDC:q <= 8'h00;
            12'h1FDD:q <= 8'h00;
            12'h1FDE:q <= 8'h00;
            12'h1FDF:q <= 8'h00;
            12'h1FE0:q <= 8'h00;
            12'h1FE1:q <= 8'h00;
            12'h1FE2:q <= 8'h00;
            12'h1FE3:q <= 8'h00;
            12'h1FE4:q <= 8'h00;
            12'h1FE5:q <= 8'h00;
            12'h1FE6:q <= 8'h00;
            12'h1FE7:q <= 8'h00;
            12'h1FE8:q <= 8'h00;
            12'h1FE9:q <= 8'h00;
            12'h1FEA:q <= 8'h00;
            12'h1FEB:q <= 8'h00;
            12'h1FEC:q <= 8'h00;
            12'h1FED:q <= 8'h00;
            12'h1FEE:q <= 8'h00;
            12'h1FEF:q <= 8'h00;
            12'h1FF0:q <= 8'h00;
            12'h1FF1:q <= 8'h00;
            12'h1FF2:q <= 8'h00;
            12'h1FF3:q <= 8'h00;
            12'h1FF4:q <= 8'h00;
            12'h1FF5:q <= 8'h00;
            12'h1FF6:q <= 8'h00;
            12'h1FF7:q <= 8'h00;
            12'h1FF8:q <= 8'h00;
            12'h1FF9:q <= 8'h00;
            12'h1FFA:q <= 8'h00;
            12'h1FFB:q <= 8'h00;
            12'h1FFC:q <= 8'h00;
            12'h1FFD:q <= 8'h00;
            12'h1FFE:q <= 8'h00;
            12'h1FFF:q <= 8'h00;
            endcase
        end
    end    
endmodule
