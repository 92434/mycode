
`timescale 1ns / 1ps
module F_normal_t10_next_Rom7(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[159:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 160'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h13: rd_q <= 160'b1001010101010110000100000011110100111111110101111111111101111110000101010111111101111000101101110101001001101110111000011111001000111000011100100101001110010110;
			5'h12: rd_q <= 160'b0001111101010000010011011111111011001111001011100011100001001110100110110000001001100101110111001110101111100010011100101101010011111100110010000010101000110011;
			5'h11: rd_q <= 160'b1101101100100110110110000101101110101111011101011100111000101101000110001001110001111100011001011100011010001100110111011000110000110010101110010000011110011111;
			5'h10: rd_q <= 160'b0110110111001110010001000000111001101110111100101100000101001111011100011101101111001001011000100011111000001101110111110111011011000000101001110110111001110101;
			5'h0f: rd_q <= 160'b1101010110100101100001100001111100011101110111010110110000011011000001000111110011111100101001111111101111110000101001001001001101101000100100110010010110111011;
			5'h0e: rd_q <= 160'b1011010111001100100110011000100000110110111110000001001011000000001000010100001000101011101001110001000001000101001101010000100110111000000010100010100000010010;
			5'h0d: rd_q <= 160'b1110010100010101001111101110100000000110101011100100111001110011101100111000100111011101010111111010100111100110110110100000100110001101011100110001010000001100;
			5'h0c: rd_q <= 160'b1001010010100000010010001011100111101100110100001101100000100111100010010100110100100101010101101010000000110110100111111000000001001110100100010100000111010010;
			5'h0b: rd_q <= 160'b0010100001000001111000011010101001110111110100101010100010110101011101001011111011000011001011001101110011111100110101111000001101101000001011010111001101100000;
			5'h0a: rd_q <= 160'b1110111100110100010001010011010110001010111000000011111001011001011001011101000100101000001010110001011001000101100101111111100000000010000011001111101101110111;
			5'h09: rd_q <= 160'b1110110011000110111001100101111101011000000111111001011111110111101110010100001000111011100001011110011110011101100001110100000011111000110101000111100100001111;
			5'h08: rd_q <= 160'b0011100000011110000100010001110100011010011111110111111110010011101100110001001001011011110001000111110101010011011011101011010000100001000100110100001000001000;
			5'h07: rd_q <= 160'b1110011110111110011101110001010011100101100000011101101100110001001111110001100000100101010101101001000101101000111111010000001011001110001101101100111111000110;
			5'h06: rd_q <= 160'b1000011110110000101000110010011111010110001010000111010011100011111011001101111101011111000111010010110111110100101010100111000001001101111010001101001110101001;
			5'h05: rd_q <= 160'b0101000000111110011111101101110010000000101010110101000110111001101010100000001000010111011100001010010001100101101011100011101111011111111001000100110111000000;
			5'h04: rd_q <= 160'b1100110100100101100011011110110110011100001001100110010101011101100110010011010100010011011010101111010000001110000110111000111001010111011101110001100001001000;
			5'h03: rd_q <= 160'b1010001110011000001000100000011011010101011001011100011111010000000100010100011100001101001101010100001110000111100010100110100000101111110110001111111110011111;
			5'h02: rd_q <= 160'b0110110110110110111110101111010000110011100010001101000101000110100011001101001000010010000100110110111010001000110101000010000100100100101110100000111110001101;
			5'h01: rd_q <= 160'b1000100011011000001001100101110101001111111101101000101000110001011010011110011100011000011110000100011001010011010001000100001111101001011110100111001101011001;
			5'h00: rd_q <= 160'b1110101011001010101001111010000010101010110111111011011100110011101100000100101011110101001111100101100011101000110000100110001001000000010110100100100001100111;
		default:rd_q <= 160'b0;
		endcase
	end
end

endmodule
