`timescale 1ns / 1ps
module F_normal_t12_next_Rom6(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b010001111101101110111101001011010011100101111100000100000111011101100111100110010011010101100000000101101000100011011001101110110001100100001101000110001101001000001011111101101110110011110011;
			5'h16: rd_q <= 192'b101001101100010000100000011101010000000101000110110000100111010000000100010001001010010001010111110000110100010101101100000101101101111100101011011010100100111001010101000001000001110110000110;
			5'h15: rd_q <= 192'b001011110110000001000011001100011101000100100100100101001001101101001101101111111011011100111111011101110110111011011100101010110000010101000010001110000011110110010011001111100101010101111010;
			5'h14: rd_q <= 192'b010101010111101100110001011001001011101110100011000101101001011111100111111001111001010110010011111110110010101001100110001101100101011010010001101111100000110000010010010111001101100001101111;
			5'h13: rd_q <= 192'b011100011101000110100110100000110100010100001010100101100011100001011100000010011101001001100000100001000011101111101001110010010001011010000000101100000011001000101000001011010100111110111000;
			5'h12: rd_q <= 192'b100001101000000101011101111110011010100000111010001110110100001011111010111101111110110010110000001001001111111101100000001101110000100101000000010000110110011100110111110110010111000111001101;
			5'h11: rd_q <= 192'b000011110011001101110001110110110101101010001101011001111101001011001010110010011101110001110111011101111010000111011001101101101000000011110000111101111001010100111000101000100011111111111110;
			5'h10: rd_q <= 192'b001111010100011001011000011010101100110001110001011111010100101011110000010000100010010100000011100001010000111111101001010011110100000110000100000001110100011001101100011010101111100110010001;
			5'h0f: rd_q <= 192'b010011001111000011110000111100010101110001010110101101000111111010100011100101101001101100001111111001100011110110000100110100001001100010010011010100100011101010011011000000010010001000110111;
			5'h0e: rd_q <= 192'b101111010000011100010001001101110011011110101010110110111001111000011011001010100011101100011111000101110000101011100000101100101010001001111111111000101001000110001011101100010110010111100101;
			5'h0d: rd_q <= 192'b000000010111001001010011100100011111101011101000111010010001111000011111001110010000101101100011011010010010000101100011000001101010011011010011011010111001011011010010000010010101000110101101;
			5'h0c: rd_q <= 192'b101000100010000101110010100110010001000101000110110111100001000001101011111100001100001110111000111101001000111110110001111110000001101110110010110011010000010010011000110100111010000010001001;
			5'h0b: rd_q <= 192'b111100110111010110001011100111010011111100011100110010101011100100011111111000101110011110000101110111111111101001100011100101000110000110111101001010011010111110101100010110001101111011110000;
			5'h0a: rd_q <= 192'b001001011110110010101101100111101111101100100011010110000010001010001111011110011101110001101110001000000111010001011000110000000101110101010010011101001110010111100111110111100100110101001100;
			5'h09: rd_q <= 192'b001011000111110111000010101111011010000101100000011101101000101000011001011100001100100011110111101000101110000100111110010100111111101100100010011010011100101110111111100010010100111010111011;
			5'h08: rd_q <= 192'b000001010100000011010010010000001101110010111101101010110010111000001101111101111001011001000001101101010010000111111100100011000011111010101100010011110010010000000001001100110010101100110100;
			5'h07: rd_q <= 192'b001111101101001010000010110010001100110001001001110010100000110100001110110000010101100111111001010111111010000110111010101001100101001111011000011100110001011001011010010101101010100100010100;
			5'h06: rd_q <= 192'b111000001010100111000000111001110001000000010000101001000001110010011000100101101110100000000011001110101011001011110101001010001100111100011101101100111000001111011001001000011011000111111000;
			5'h05: rd_q <= 192'b111101011100010100000101101011001011101110111111110100000001000010010110101110110010010110010111110010101101101110010000101011101111010011011100110000110111010001100110100100000100111100001010;
			5'h04: rd_q <= 192'b100101110001010000001100010100011010111101110100001010111111101111001011010010100000001110110011111011010000100010000010110100111010001011011001110100110001101011010010101010110000011110010101;
			5'h03: rd_q <= 192'b110000111110110111011000111111110001010111001101100100011100011011011101100111111111100111101001011110110100010000110000110011010011011001101010001111100100101011010000010100100011101000101111;
			5'h02: rd_q <= 192'b000000101001001000010000010110011010100101110100000010011101111101000101101110111111110000010001011100110010000111111110000110101111000110100101010101101010001010001110010101110111001101100011;
			5'h01: rd_q <= 192'b001011100000101101000001100000010011000001010011111001011001010101100111110111000110100100111111010001111110100011010001110111110001110100011101101000100111010100111100011001111110011011011100;
			5'h00: rd_q <= 192'b101001001111110000001101000010001111101100101110001010011100111101100101001000101000001011100011000001100100111010110110001101001000011110111100010001100110100000110110101101001010110111010101;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
