`timescale 1ns / 1ps
module F_normal_t12_next_Rom5(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b100011111011011101111010010110100111001011111000001000001110111011001111001100100110101011000000001011010001000110110011011101100011001000011010001100011010010000010111111011011101100111100110;
			5'h16: rd_q <= 192'b100000101101110011000000001001111101110111001110010000010110100100101010101010000001000011011001101100001110001100111110001110011100111101000010101000001101111100101000111010001111001111101001;
			5'h15: rd_q <= 192'b010111101100000010000110011000111010001001001001001010010011011010011011011111110110111001111110111011101101110110111001010101100000101010000100011100000111101100100110011111001010101011110100;
			5'h14: rd_q <= 192'b101010101111011001100010110010010111011101000110001011010010111111001111110011110010101100100111111101100101010011001100011011001010110100100011011111000001100000100100101110011011000011011110;
			5'h13: rd_q <= 192'b111000111010001101001101000001101000101000010101001011000111000010111000000100111010010011000001000010000111011111010011100100100010110100000001011000000110010001010000010110101001111101110000;
			5'h12: rd_q <= 192'b110000100101011000111011001111101000111100110111101100110000010011010111110011101000000100010110011111111001011100100110011110100110001110010100111100101000110111101101010100100010101101111111;
			5'h11: rd_q <= 192'b000111100110011011100011101101101011010100011010110011111010010110010101100100111011100011101110111011110100001110110011011011010000000111100001111011110010101001110001010001000111111111111100;
			5'h10: rd_q <= 192'b011110101000110010110000110101011001100011100010111110101001010111100000100001000100101000000111000010100001111111010010100111101000001100001000000011101000110011011000110101011111001100100010;
			5'h0f: rd_q <= 192'b100110011110000111100001111000101011100010101101011010001111110101000111001011010011011000011111110011000111101100001001101000010011000100100110101001000111010100110110000000100100010001101110;
			5'h0e: rd_q <= 192'b101101010101101010100010101000111011000000010110011100101011110100010100011101010010111001001000000110000111110000100111011100010011010111101011101100010110000010010101100000100000001100101111;
			5'h0d: rd_q <= 192'b000000101110010010100111001000111111010111010001110100100011110000111110011100100001011011000110110100100100001011000110000011010100110110100110110101110010110110100100000100101010001101011010;
			5'h0c: rd_q <= 192'b100010110001011001100101111111111111110111001110011110011010000111110101110000001101111100000111110111110111011010000101111001000100011001110001111011100100101010110011010001111000100111110111;
			5'h0b: rd_q <= 192'b001010011011111110010111111101111010000101111010010100001111001100011101111001001001011101111101100010011001110100100001001111001011001001101110001001110001110011011010010100010111010100000101;
			5'h0a: rd_q <= 192'b010010111101100101011011001111011111011001000110101100000100010100011110111100111011100011011100010000001110100010110001100000001011101010100100111010011100101111001111101111001001101010011000;
			5'h09: rd_q <= 192'b010110001111101110000101011110110100001011000000111011010001010000110010111000011001000111101111010001011100001001111100101001111111011001000100110100111001011101111111000100101001110101110110;
			5'h08: rd_q <= 192'b000010101000000110100100100000011011100101111011010101100101110000011011111011110010110010000011011010100100001111111001000110000111110101011000100111100100100000000010011001100101011001101000;
			5'h07: rd_q <= 192'b011111011010010100000101100100011001100010010011100101000001101000011101100000101011001111110010101111110100001101110101010011001010011110110000111001100010110010110100101011010101001000101000;
			5'h06: rd_q <= 192'b000011100000011100000001000000111111111101100010100011011011100000010011000011001000100001110000010000110000110000001100010001011110111100101111000100110100010000110000101000111010101100010101;
			5'h05: rd_q <= 192'b001001001101111010001011100101001010100000111100011001011010000000001111010101110001001101011001101000111101111011000111010010011001100010101101111100101010101101001111110000000101011011110001;
			5'h04: rd_q <= 192'b111000010111110010011000011011101000000110101011100100100111011010110100101101010101111100010001111011000111100011100011101100110011010010100111110100100111011000100111101101101100011111001111;
			5'h03: rd_q <= 192'b010010001000111100110001001100111111010011011000111001100000110010011001000111101010101110100100110000001110000110000111100011100001110111000000000010001101011000100010010001001011110010111011;
			5'h02: rd_q <= 192'b000001010010010000100000101100110101001011101000000100111011111010001011011101111111100000100010111001100100001111111100001101011110001101001010101011010100010100011100101011101110011011000110;
			5'h01: rd_q <= 192'b010111000001011010000011000000100110000010100111110010110010101011001111101110001101001001111110100011111101000110100011101111100011101000111011010001001110101001111000110011111100110110111000;
			5'h00: rd_q <= 192'b100001101010110010011010110111000010100100011111100101100001111111101000011001000101110110110000001110101111010010001010011111010111111001101100111110001001001111101111100010011001001101001111;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
