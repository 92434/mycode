`timescale 1 ns / 1 ps

module ck_processer #(
		parameter integer AXI_DATA_WIDTH = 32,
		parameter integer CSA_CALC_IN_WIDTH = 8 * 8,
		parameter integer CYPHER_DATA_WIDTH = 8 * 8
	)
	(
		input wire init,
		input wire [31 : 0] block,
		input wire [CSA_CALC_IN_WIDTH - 1 : 0] in,
		input wire [CYPHER_DATA_WIDTH - 1 : 0] cb,
		input wire [AXI_DATA_WIDTH - 1 : 0] loops,

		output wire [CYPHER_DATA_WIDTH - 1 : 0] ck_out
	);
	reg[2047:0] box={
		8'h22,
		8'hcc,
		8'he3,
		8'hbd,
		8'h36,
		8'h8a,
		8'hde,
		8'h65,
		8'h1a,
		8'hd9,
		8'h3f,
		8'h10,
		8'h20,
		8'h0b,
		8'h80,
		8'hbf,
		8'h21,
		8'h04,
		8'h54,
		8'h32,
		8'ha9,
		8'h3d,
		8'h90,
		8'h38,
		8'hcd,
		8'h1c,
		8'h66,
		8'had,
		8'h85,
		8'h72,
		8'hd8,
		8'hc1,
		8'hc7,
		8'h1d,
		8'h9a,
		8'h29,
		8'h5b,
		8'h4e,
		8'h5d,
		8'h7d,
		8'h8d,
		8'hdc,
		8'hb8,
		8'hf3,
		8'h50,
		8'h8b,
		8'hf4,
		8'h9e,
		8'h62,
		8'h8e,
		8'h23,
		8'hfd,
		8'h30,
		8'h06,
		8'h7e,
		8'h99,
		8'h69,
		8'hf8,
		8'h5e,
		8'h46,
		8'hd4,
		8'ha3,
		8'he0,
		8'hce,
		8'hc3,
		8'hf5,
		8'h0e,
		8'hfe,
		8'hcb,
		8'h2a,
		8'hac,
		8'hb0,
		8'h8f,
		8'hbc,
		8'heb,
		8'hca,
		8'h88,
		8'h0a,
		8'ha2,
		8'hab,
		8'hee,
		8'hd5,
		8'hef,
		8'h91,
		8'h5c,
		8'h9c,
		8'hf9,
		8'haf,
		8'hb2,
		8'h2f,
		8'h61,
		8'hff,
		8'h35,
		8'h2d,
		8'hc8,
		8'h86,
		8'h4d,
		8'h53,
		8'hbb,
		8'h00,
		8'hba,
		8'ha0,
		8'hb4,
		8'h92,
		8'hed,
		8'h9b,
		8'h97,
		8'h7f,
		8'he8,
		8'h4a,
		8'h63,
		8'h6d,
		8'he2,
		8'hda,
		8'hdf,
		8'hf2,
		8'ha5,
		8'h98,
		8'hb3,
		8'hd2,
		8'h40,
		8'hc6,
		8'h3a,
		8'ha7,
		8'h70,
		8'hf7,
		8'h79,
		8'hf6,
		8'h48,
		8'h3c,
		8'h0f,
		8'h71,
		8'h68,
		8'h82,
		8'h95,
		8'hd6,
		8'h76,
		8'h09,
		8'h18,
		8'h03,
		8'hae,
		8'h31,
		8'h67,
		8'h33,
		8'h7c,
		8'hdd,
		8'h45,
		8'h93,
		8'hf0,
		8'hd3,
		8'h6a,
		8'h58,
		8'h57,
		8'hc4,
		8'h52,
		8'he5,
		8'h73,
		8'hf1,
		8'hcf,
		8'h94,
		8'hd1,
		8'ha6,
		8'h78,
		8'h41,
		8'h83,
		8'h0d,
		8'h51,
		8'hdb,
		8'h5f,
		8'hc9,
		8'h14,
		8'h7b,
		8'hd0,
		8'h0c,
		8'h77,
		8'hb9,
		8'hea,
		8'h12,
		8'h19,
		8'hc2,
		8'h55,
		8'h17,
		8'he6,
		8'h64,
		8'h9f,
		8'h1e,
		8'hb1,
		8'hfa,
		8'h1b,
		8'hd7,
		8'he4,
		8'h59,
		8'h49,
		8'h37,
		8'h28,
		8'haa,
		8'h11,
		8'hc5,
		8'h60,
		8'hb6,
		8'h6c,
		8'h75,
		8'h02,
		8'h2c,
		8'h43,
		8'h47,
		8'hec,
		8'hbe,
		8'hfc,
		8'h01,
		8'h6f,
		8'h1f,
		8'h08,
		8'ha4,
		8'h05,
		8'ha8,
		8'h44,
		8'h26,
		8'he1,
		8'h07,
		8'h84,
		8'hb5,
		8'h6e,
		8'h8c,
		8'h2b,
		8'h25,
		8'h42,
		8'h87,
		8'h6b,
		8'h7a,
		8'h89,
		8'h9d,
		8'h4b,
		8'h74,
		8'h16,
		8'ha1,
		8'h3e,
		8'h24,
		8'h13,
		8'hfb,
		8'he7,
		8'h81,
		8'h2e,
		8'hc0,
		8'h3b,
		8'h4f,
		8'h4c,
		8'h15,
		8'h56,
		8'h27,
		8'h96,
		8'h5a,
		8'hb7,
		8'h34,
		8'he9,
		8'h39
	};
	
	assign ck_out[7:0]  =(init==1)?in[7:0]:(((block[31:30]==2'b01)?(box[((in[7:0]+in[55:48])%256)*8+:8]^in[7:0]):(box[((cb[7:0]+cb[55:48])%256)*8+:8]^cb[7:0]))^(loops));
	assign ck_out[15:8] =(init==1)?in[15:8]:(((block[31:30]==2'b01)?(box[((in[15:8]+in[55:48])%256)*8+:8]^in[15:8]):(box[((cb[15:8]+cb[55:48])%256)*8+:8]^cb[15:8]))^(loops>>8));
	assign ck_out[23:16]=(init==1)?in[23:16]:((block[31:30]==2'b01)?(box[((in[23:16]+in[55:48])%256)*8+:8]^in[23:16]):(box[((cb[23:16]+cb[55:48])%256)*8+:8]^cb[23:16]));
	assign ck_out[31:24]=(init==1)?in[7:0]+in[15:8]+in[23:16]:((block[31:30]==2'b01)?(((box[((in[7:0]+in[55:48])%256)*8+:8]^in[7:0])^loops)+((box[((in[15:8]+in[55:48])%256)*8+:8]^in[15:8])^(loops>>8))+(box[((in[23:16]+in[55:48])%256)*8+:8]^in[23:16])):(((box[((cb[7:0]+cb[55:48])%256)*8+:8]^cb[7:0])^loops)+((box[((cb[15:8]+cb[55:48])%256)*8+:8]^cb[15:8])^(loops>>8))+(box[((cb[23:16]+cb[55:48])%256)*8+:8]^cb[23:16])));
	assign ck_out[39:32]=(init==1)?in[31:24]:((block[31:30]==2'b01)?(box[((in[31:24]+in[55:48])%256)*8+:8]^in[31:24]):(box[((cb[31:24]+cb[55:48])%256)*8+:8]^cb[31:24]));
	assign ck_out[47:40]=(init==1)?in[39:32]:((block[31:30]==2'b01)?(box[((in[39:32]+in[55:48])%256)*8+:8]^in[39:32]):(box[((cb[39:32]+cb[55:48])%256)*8+:8]^cb[39:32]));
	assign ck_out[55:48]=(init==1)?0:((block[31:30]==2'b01)?(box[((in[47:40]+in[55:48])%256)*8+:8]^in[47:40]):(box[((cb[47:40]+cb[55:48])%256)*8+:8]^cb[47:40]));
	assign ck_out[63:56]=(init==1)?in[31:24]+in[39:32]:((block[31:30]==2'b01)?((box[((in[31:24]+in[55:48])%256)*8+:8]^in[31:24])+(box[((in[39:32]+in[55:48])%256)*8+:8]^in[39:32])+(box[((in[47:40]+in[55:48])%256)*8+:8]^in[47:40])):((box[((cb[31:24]+cb[55:48])%256)*8+:8]^cb[31:24])+(box[((cb[39:32]+cb[55:48])%256)*8+:8]^cb[39:32])+(box[((cb[47:40]+cb[55:48])%256)*8+:8]^cb[47:40])));

endmodule
