
`timescale 1ns / 1ps
module F_normal_t8_next_Rom5(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[127:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 128'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h0f: rd_q <= 128'b10111000111101101110010001001001111111001001100010010001101010000010011011110010010110011110110111110000001000111011011100100101;
			5'h0e: rd_q <= 128'b11001001010110010100001111100111101101101011010010111101011110011111011011100110101101101010101110100010001000000011000101001001;
			5'h0d: rd_q <= 128'b11110111110101000001011010000011001111001100110111001100101101100100011001111101000010100000101111000010101001000110001111000011;
			5'h0c: rd_q <= 128'b01110010101100010001111100100000000000100101011010100001011100101010110010000011110001111000011110001111110110111001001000111000;
			5'h0b: rd_q <= 128'b11110110110001110011001111100001101110100010010001000010110101010111110001011100101111001011001111110011011111001101000110100000;
			5'h0a: rd_q <= 128'b11100001100010011111111111011011011001001010000110010100001111000100011111101111110000010001000111110111111111101010010011100111;
			5'h09: rd_q <= 128'b11111111010010000000000101001000100011010011101111010011011001000010111100001010011101011000001011011011011001000100011111010100;
			5'h08: rd_q <= 128'b00011100110100001010111100011100010110000010111001001101110111001011011001111101011110011100000000101010010110101101111101000001;
			5'h07: rd_q <= 128'b00101110001000010110100110111101011000110111111000001010001001111101010100001010111010110000001010111100001000101011011100010110;
			5'h06: rd_q <= 128'b00101010010010011111101111000000000001001101011101011111000111011011100000001010101001111110111100101111011111100011001000111111;
			5'h05: rd_q <= 128'b10000010011110100011010011001010110111100011110100011110011010011100110001100010110000000111101001101000000100000110010101011010;
			5'h04: rd_q <= 128'b00100001000000001111110110010110011111001111010011001110000011001011100000100010000111101010100011001111110101010110100111101111;
			5'h03: rd_q <= 128'b00100110101010000111111010011000011001000111111011011010010111110010100111000010110000101001101101110111010100101100001000100010;
			5'h02: rd_q <= 128'b10111101001000101110001010110010111000110011001110000110011100001101111011000011011100111001100100100111011010110101000101100110;
			5'h01: rd_q <= 128'b01101111011111001100001111110111011000100111011101000101010010001000100100110010110110011000001010101000010010101010111111001100;
			5'h00: rd_q <= 128'b11011111111011001011111011101000010101100100101010011010110110001011101101010001000001110011101111100000011100111100001110010101;
		default:rd_q <= 128'b0;
		endcase
	end
end

endmodule
