
`timescale 1ns / 1ps
module order_ctrl(
input	          							sys_clk,
input											fs_en,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input	          							frame_mode,
input	          			[3:0] 		ldpc_mode,
input	          			[2:0] 		order_idx,
input	          							shift_vld,
//////////////////////////////////////////////////////////////
input	          			[359:0] 		order_in,
output      reg   		[359:0] 		order_out
);

reg 							[2:0]			mode_switch_tmp;

always @(posedge sys_clk)begin
	if(~rst_n)begin
		mode_switch_tmp <= 3'b000;
	end
	else begin
	case({ldpc_mode,frame_mode})
		5'b00000:mode_switch_tmp <= 3'b000;//00 51
		5'b01011:mode_switch_tmp <= 3'b000;
		5'b00101:mode_switch_tmp <= 3'b001;//21
		5'b00111:mode_switch_tmp <= 3'b010;//31
		5'b01100:mode_switch_tmp <= 3'b011;//60 91
		5'b10011:mode_switch_tmp <= 3'b011;
		5'b00001:mode_switch_tmp <= 3'b100;//01 20 50 61 70 90
		5'b00100:mode_switch_tmp <= 3'b100;
		5'b01010:mode_switch_tmp <= 3'b100;
		5'b01101:mode_switch_tmp <= 3'b100;
		5'b01110:mode_switch_tmp <= 3'b100;
		5'b10010:mode_switch_tmp <= 3'b100;
		5'b00010:mode_switch_tmp <= 3'b101;//10 40 81
		5'b01000:mode_switch_tmp <= 3'b101;
		5'b10001:mode_switch_tmp <= 3'b101;
		5'b00011:mode_switch_tmp <= 3'b110;//11 80
		5'b10000:mode_switch_tmp <= 3'b110;
		5'b00110:mode_switch_tmp <= 3'b111;//30 41 71 100
		5'b01001:mode_switch_tmp <= 3'b111;
		5'b01111:mode_switch_tmp <= 3'b111;
		5'b10100:mode_switch_tmp <= 3'b111;
		default:mode_switch_tmp <= 3'b000;
	endcase
	end
end

always @(posedge sys_clk)begin
	if(~rst_n)begin
		order_out <= 360'h00;
	end
	else if(fs_en == 1'b1)begin
		if(shift_vld)begin
			case({mode_switch_tmp,order_idx})
			6'b000000: order_out <= {order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6]};
			6'b000001: order_out <= {order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5]};
			6'b000010: order_out <= {order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4]};
			6'b000011: order_out <= {order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3]};
			6'b000100: order_out <= {order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2]};
			6'b000101: order_out <= {order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1]};
			6'b000110: order_out <= {order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0]};
			6'b000111: order_out <= {order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7]};
			6'b001000: order_out <= {order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2]};
			6'b001001: order_out <= {order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5]};
			6'b001010: order_out <= {order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0]};
			6'b001011: order_out <= {order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3]};
			6'b001100: order_out <= {order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6]};
			6'b001101: order_out <= {order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1]};
			6'b001110: order_out <= {order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4]};
			6'b001111: order_out <= {order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7]};
			6'b010000: order_out <= {order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0]};
			6'b010001: order_out <= {order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1]};
			6'b010010: order_out <= {order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2]};
			6'b010011: order_out <= {order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3]};
			6'b010100: order_out <= {order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4]};
			6'b010101: order_out <= {order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5]};
			6'b010110: order_out <= {order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6]};
			6'b010111: order_out <= {order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7]};
			6'b011000: order_out <= {order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4]};
			6'b011001: order_out <= {order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1]};
			6'b011010: order_out <= {order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6]};
			6'b011011: order_out <= {order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3]};
			6'b011100: order_out <= {order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0]};
			6'b011101: order_out <= {order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5]};
			6'b011110: order_out <= {order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7],order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2]};
			6'b011111: order_out <= {order_in[354],order_in[346],order_in[338],order_in[330],order_in[322],order_in[314],order_in[306],order_in[298],order_in[290],order_in[282],order_in[274],order_in[266],order_in[258],order_in[250],order_in[242],order_in[234],order_in[226],order_in[218],order_in[210],order_in[202],order_in[194],order_in[186],order_in[178],order_in[170],order_in[162],order_in[154],order_in[146],order_in[138],order_in[130],order_in[122],order_in[114],order_in[106],order_in[98],order_in[90],order_in[82],order_in[74],order_in[66],order_in[58],order_in[50],order_in[42],order_in[34],order_in[26],order_in[18],order_in[10],order_in[2],order_in[357],order_in[349],order_in[341],order_in[333],order_in[325],order_in[317],order_in[309],order_in[301],order_in[293],order_in[285],order_in[277],order_in[269],order_in[261],order_in[253],order_in[245],order_in[237],order_in[229],order_in[221],order_in[213],order_in[205],order_in[197],order_in[189],order_in[181],order_in[173],order_in[165],order_in[157],order_in[149],order_in[141],order_in[133],order_in[125],order_in[117],order_in[109],order_in[101],order_in[93],order_in[85],order_in[77],order_in[69],order_in[61],order_in[53],order_in[45],order_in[37],order_in[29],order_in[21],order_in[13],order_in[5],order_in[352],order_in[344],order_in[336],order_in[328],order_in[320],order_in[312],order_in[304],order_in[296],order_in[288],order_in[280],order_in[272],order_in[264],order_in[256],order_in[248],order_in[240],order_in[232],order_in[224],order_in[216],order_in[208],order_in[200],order_in[192],order_in[184],order_in[176],order_in[168],order_in[160],order_in[152],order_in[144],order_in[136],order_in[128],order_in[120],order_in[112],order_in[104],order_in[96],order_in[88],order_in[80],order_in[72],order_in[64],order_in[56],order_in[48],order_in[40],order_in[32],order_in[24],order_in[16],order_in[8],order_in[0],order_in[355],order_in[347],order_in[339],order_in[331],order_in[323],order_in[315],order_in[307],order_in[299],order_in[291],order_in[283],order_in[275],order_in[267],order_in[259],order_in[251],order_in[243],order_in[235],order_in[227],order_in[219],order_in[211],order_in[203],order_in[195],order_in[187],order_in[179],order_in[171],order_in[163],order_in[155],order_in[147],order_in[139],order_in[131],order_in[123],order_in[115],order_in[107],order_in[99],order_in[91],order_in[83],order_in[75],order_in[67],order_in[59],order_in[51],order_in[43],order_in[35],order_in[27],order_in[19],order_in[11],order_in[3],order_in[358],order_in[350],order_in[342],order_in[334],order_in[326],order_in[318],order_in[310],order_in[302],order_in[294],order_in[286],order_in[278],order_in[270],order_in[262],order_in[254],order_in[246],order_in[238],order_in[230],order_in[222],order_in[214],order_in[206],order_in[198],order_in[190],order_in[182],order_in[174],order_in[166],order_in[158],order_in[150],order_in[142],order_in[134],order_in[126],order_in[118],order_in[110],order_in[102],order_in[94],order_in[86],order_in[78],order_in[70],order_in[62],order_in[54],order_in[46],order_in[38],order_in[30],order_in[22],order_in[14],order_in[6],order_in[353],order_in[345],order_in[337],order_in[329],order_in[321],order_in[313],order_in[305],order_in[297],order_in[289],order_in[281],order_in[273],order_in[265],order_in[257],order_in[249],order_in[241],order_in[233],order_in[225],order_in[217],order_in[209],order_in[201],order_in[193],order_in[185],order_in[177],order_in[169],order_in[161],order_in[153],order_in[145],order_in[137],order_in[129],order_in[121],order_in[113],order_in[105],order_in[97],order_in[89],order_in[81],order_in[73],order_in[65],order_in[57],order_in[49],order_in[41],order_in[33],order_in[25],order_in[17],order_in[9],order_in[1],order_in[356],order_in[348],order_in[340],order_in[332],order_in[324],order_in[316],order_in[308],order_in[300],order_in[292],order_in[284],order_in[276],order_in[268],order_in[260],order_in[252],order_in[244],order_in[236],order_in[228],order_in[220],order_in[212],order_in[204],order_in[196],order_in[188],order_in[180],order_in[172],order_in[164],order_in[156],order_in[148],order_in[140],order_in[132],order_in[124],order_in[116],order_in[108],order_in[100],order_in[92],order_in[84],order_in[76],order_in[68],order_in[60],order_in[52],order_in[44],order_in[36],order_in[28],order_in[20],order_in[12],order_in[4],order_in[359],order_in[351],order_in[343],order_in[335],order_in[327],order_in[319],order_in[311],order_in[303],order_in[295],order_in[287],order_in[279],order_in[271],order_in[263],order_in[255],order_in[247],order_in[239],order_in[231],order_in[223],order_in[215],order_in[207],order_in[199],order_in[191],order_in[183],order_in[175],order_in[167],order_in[159],order_in[151],order_in[143],order_in[135],order_in[127],order_in[119],order_in[111],order_in[103],order_in[95],order_in[87],order_in[79],order_in[71],order_in[63],order_in[55],order_in[47],order_in[39],order_in[31],order_in[23],order_in[15],order_in[7]};
			6'b100000: order_out <= {order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0]};
			6'b100001: order_out <= {order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90]};
			6'b100010: order_out <= {order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180]};
			6'b100011: order_out <= {order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270]};
			6'b100100: order_out <= {order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1]};
			6'b100101: order_out <= {order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91]};
			6'b100110: order_out <= {order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271],order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181]};
			6'b100111: order_out <= {order_in[269],order_in[267],order_in[265],order_in[263],order_in[261],order_in[259],order_in[257],order_in[255],order_in[253],order_in[251],order_in[249],order_in[247],order_in[245],order_in[243],order_in[241],order_in[239],order_in[237],order_in[235],order_in[233],order_in[231],order_in[229],order_in[227],order_in[225],order_in[223],order_in[221],order_in[219],order_in[217],order_in[215],order_in[213],order_in[211],order_in[209],order_in[207],order_in[205],order_in[203],order_in[201],order_in[199],order_in[197],order_in[195],order_in[193],order_in[191],order_in[189],order_in[187],order_in[185],order_in[183],order_in[181],order_in[179],order_in[177],order_in[175],order_in[173],order_in[171],order_in[169],order_in[167],order_in[165],order_in[163],order_in[161],order_in[159],order_in[157],order_in[155],order_in[153],order_in[151],order_in[149],order_in[147],order_in[145],order_in[143],order_in[141],order_in[139],order_in[137],order_in[135],order_in[133],order_in[131],order_in[129],order_in[127],order_in[125],order_in[123],order_in[121],order_in[119],order_in[117],order_in[115],order_in[113],order_in[111],order_in[109],order_in[107],order_in[105],order_in[103],order_in[101],order_in[99],order_in[97],order_in[95],order_in[93],order_in[91],order_in[89],order_in[87],order_in[85],order_in[83],order_in[81],order_in[79],order_in[77],order_in[75],order_in[73],order_in[71],order_in[69],order_in[67],order_in[65],order_in[63],order_in[61],order_in[59],order_in[57],order_in[55],order_in[53],order_in[51],order_in[49],order_in[47],order_in[45],order_in[43],order_in[41],order_in[39],order_in[37],order_in[35],order_in[33],order_in[31],order_in[29],order_in[27],order_in[25],order_in[23],order_in[21],order_in[19],order_in[17],order_in[15],order_in[13],order_in[11],order_in[9],order_in[7],order_in[5],order_in[3],order_in[1],order_in[358],order_in[356],order_in[354],order_in[352],order_in[350],order_in[348],order_in[346],order_in[344],order_in[342],order_in[340],order_in[338],order_in[336],order_in[334],order_in[332],order_in[330],order_in[328],order_in[326],order_in[324],order_in[322],order_in[320],order_in[318],order_in[316],order_in[314],order_in[312],order_in[310],order_in[308],order_in[306],order_in[304],order_in[302],order_in[300],order_in[298],order_in[296],order_in[294],order_in[292],order_in[290],order_in[288],order_in[286],order_in[284],order_in[282],order_in[280],order_in[278],order_in[276],order_in[274],order_in[272],order_in[270],order_in[268],order_in[266],order_in[264],order_in[262],order_in[260],order_in[258],order_in[256],order_in[254],order_in[252],order_in[250],order_in[248],order_in[246],order_in[244],order_in[242],order_in[240],order_in[238],order_in[236],order_in[234],order_in[232],order_in[230],order_in[228],order_in[226],order_in[224],order_in[222],order_in[220],order_in[218],order_in[216],order_in[214],order_in[212],order_in[210],order_in[208],order_in[206],order_in[204],order_in[202],order_in[200],order_in[198],order_in[196],order_in[194],order_in[192],order_in[190],order_in[188],order_in[186],order_in[184],order_in[182],order_in[180],order_in[178],order_in[176],order_in[174],order_in[172],order_in[170],order_in[168],order_in[166],order_in[164],order_in[162],order_in[160],order_in[158],order_in[156],order_in[154],order_in[152],order_in[150],order_in[148],order_in[146],order_in[144],order_in[142],order_in[140],order_in[138],order_in[136],order_in[134],order_in[132],order_in[130],order_in[128],order_in[126],order_in[124],order_in[122],order_in[120],order_in[118],order_in[116],order_in[114],order_in[112],order_in[110],order_in[108],order_in[106],order_in[104],order_in[102],order_in[100],order_in[98],order_in[96],order_in[94],order_in[92],order_in[90],order_in[88],order_in[86],order_in[84],order_in[82],order_in[80],order_in[78],order_in[76],order_in[74],order_in[72],order_in[70],order_in[68],order_in[66],order_in[64],order_in[62],order_in[60],order_in[58],order_in[56],order_in[54],order_in[52],order_in[50],order_in[48],order_in[46],order_in[44],order_in[42],order_in[40],order_in[38],order_in[36],order_in[34],order_in[32],order_in[30],order_in[28],order_in[26],order_in[24],order_in[22],order_in[20],order_in[18],order_in[16],order_in[14],order_in[12],order_in[10],order_in[8],order_in[6],order_in[4],order_in[2],order_in[0],order_in[359],order_in[357],order_in[355],order_in[353],order_in[351],order_in[349],order_in[347],order_in[345],order_in[343],order_in[341],order_in[339],order_in[337],order_in[335],order_in[333],order_in[331],order_in[329],order_in[327],order_in[325],order_in[323],order_in[321],order_in[319],order_in[317],order_in[315],order_in[313],order_in[311],order_in[309],order_in[307],order_in[305],order_in[303],order_in[301],order_in[299],order_in[297],order_in[295],order_in[293],order_in[291],order_in[289],order_in[287],order_in[285],order_in[283],order_in[281],order_in[279],order_in[277],order_in[275],order_in[273],order_in[271]};
			6'b101000: order_out <= {order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0]};
			6'b101001: order_out <= {order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45]};
			6'b101010: order_out <= {order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90]};
			6'b101011: order_out <= {order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135]};
			6'b101100: order_out <= {order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180]};
			6'b101101: order_out <= {order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225]};
			6'b101110: order_out <= {order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315],order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270]};
			6'b101111: order_out <= {order_in[314],order_in[313],order_in[312],order_in[311],order_in[310],order_in[309],order_in[308],order_in[307],order_in[306],order_in[305],order_in[304],order_in[303],order_in[302],order_in[301],order_in[300],order_in[299],order_in[298],order_in[297],order_in[296],order_in[295],order_in[294],order_in[293],order_in[292],order_in[291],order_in[290],order_in[289],order_in[288],order_in[287],order_in[286],order_in[285],order_in[284],order_in[283],order_in[282],order_in[281],order_in[280],order_in[279],order_in[278],order_in[277],order_in[276],order_in[275],order_in[274],order_in[273],order_in[272],order_in[271],order_in[270],order_in[269],order_in[268],order_in[267],order_in[266],order_in[265],order_in[264],order_in[263],order_in[262],order_in[261],order_in[260],order_in[259],order_in[258],order_in[257],order_in[256],order_in[255],order_in[254],order_in[253],order_in[252],order_in[251],order_in[250],order_in[249],order_in[248],order_in[247],order_in[246],order_in[245],order_in[244],order_in[243],order_in[242],order_in[241],order_in[240],order_in[239],order_in[238],order_in[237],order_in[236],order_in[235],order_in[234],order_in[233],order_in[232],order_in[231],order_in[230],order_in[229],order_in[228],order_in[227],order_in[226],order_in[225],order_in[224],order_in[223],order_in[222],order_in[221],order_in[220],order_in[219],order_in[218],order_in[217],order_in[216],order_in[215],order_in[214],order_in[213],order_in[212],order_in[211],order_in[210],order_in[209],order_in[208],order_in[207],order_in[206],order_in[205],order_in[204],order_in[203],order_in[202],order_in[201],order_in[200],order_in[199],order_in[198],order_in[197],order_in[196],order_in[195],order_in[194],order_in[193],order_in[192],order_in[191],order_in[190],order_in[189],order_in[188],order_in[187],order_in[186],order_in[185],order_in[184],order_in[183],order_in[182],order_in[181],order_in[180],order_in[179],order_in[178],order_in[177],order_in[176],order_in[175],order_in[174],order_in[173],order_in[172],order_in[171],order_in[170],order_in[169],order_in[168],order_in[167],order_in[166],order_in[165],order_in[164],order_in[163],order_in[162],order_in[161],order_in[160],order_in[159],order_in[158],order_in[157],order_in[156],order_in[155],order_in[154],order_in[153],order_in[152],order_in[151],order_in[150],order_in[149],order_in[148],order_in[147],order_in[146],order_in[145],order_in[144],order_in[143],order_in[142],order_in[141],order_in[140],order_in[139],order_in[138],order_in[137],order_in[136],order_in[135],order_in[134],order_in[133],order_in[132],order_in[131],order_in[130],order_in[129],order_in[128],order_in[127],order_in[126],order_in[125],order_in[124],order_in[123],order_in[122],order_in[121],order_in[120],order_in[119],order_in[118],order_in[117],order_in[116],order_in[115],order_in[114],order_in[113],order_in[112],order_in[111],order_in[110],order_in[109],order_in[108],order_in[107],order_in[106],order_in[105],order_in[104],order_in[103],order_in[102],order_in[101],order_in[100],order_in[99],order_in[98],order_in[97],order_in[96],order_in[95],order_in[94],order_in[93],order_in[92],order_in[91],order_in[90],order_in[89],order_in[88],order_in[87],order_in[86],order_in[85],order_in[84],order_in[83],order_in[82],order_in[81],order_in[80],order_in[79],order_in[78],order_in[77],order_in[76],order_in[75],order_in[74],order_in[73],order_in[72],order_in[71],order_in[70],order_in[69],order_in[68],order_in[67],order_in[66],order_in[65],order_in[64],order_in[63],order_in[62],order_in[61],order_in[60],order_in[59],order_in[58],order_in[57],order_in[56],order_in[55],order_in[54],order_in[53],order_in[52],order_in[51],order_in[50],order_in[49],order_in[48],order_in[47],order_in[46],order_in[45],order_in[44],order_in[43],order_in[42],order_in[41],order_in[40],order_in[39],order_in[38],order_in[37],order_in[36],order_in[35],order_in[34],order_in[33],order_in[32],order_in[31],order_in[30],order_in[29],order_in[28],order_in[27],order_in[26],order_in[25],order_in[24],order_in[23],order_in[22],order_in[21],order_in[20],order_in[19],order_in[18],order_in[17],order_in[16],order_in[15],order_in[14],order_in[13],order_in[12],order_in[11],order_in[10],order_in[9],order_in[8],order_in[7],order_in[6],order_in[5],order_in[4],order_in[3],order_in[2],order_in[1],order_in[0],order_in[359],order_in[358],order_in[357],order_in[356],order_in[355],order_in[354],order_in[353],order_in[352],order_in[351],order_in[350],order_in[349],order_in[348],order_in[347],order_in[346],order_in[345],order_in[344],order_in[343],order_in[342],order_in[341],order_in[340],order_in[339],order_in[338],order_in[337],order_in[336],order_in[335],order_in[334],order_in[333],order_in[332],order_in[331],order_in[330],order_in[329],order_in[328],order_in[327],order_in[326],order_in[325],order_in[324],order_in[323],order_in[322],order_in[321],order_in[320],order_in[319],order_in[318],order_in[317],order_in[316],order_in[315]};
			6'b110000: order_out <= {order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2]};
			6'b110001: order_out <= {order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182]};
			6'b110010: order_out <= {order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1]};
			6'b110011: order_out <= {order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181]};
			6'b110100: order_out <= {order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0]};
			6'b110101: order_out <= {order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180]};
			6'b110110: order_out <= {order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3]};
			6'b110111: order_out <= {order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183]};
			6'b111000: order_out <= {order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0]};
			6'b111001: order_out <= {order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180]};
			6'b111010: order_out <= {order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1]};
			6'b111011: order_out <= {order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181]};
			6'b111100: order_out <= {order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2]};
			6'b111101: order_out <= {order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182]};
			6'b111110: order_out <= {order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183],order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3]};
			6'b111111: order_out <= {order_in[179],order_in[175],order_in[171],order_in[167],order_in[163],order_in[159],order_in[155],order_in[151],order_in[147],order_in[143],order_in[139],order_in[135],order_in[131],order_in[127],order_in[123],order_in[119],order_in[115],order_in[111],order_in[107],order_in[103],order_in[99],order_in[95],order_in[91],order_in[87],order_in[83],order_in[79],order_in[75],order_in[71],order_in[67],order_in[63],order_in[59],order_in[55],order_in[51],order_in[47],order_in[43],order_in[39],order_in[35],order_in[31],order_in[27],order_in[23],order_in[19],order_in[15],order_in[11],order_in[7],order_in[3],order_in[358],order_in[354],order_in[350],order_in[346],order_in[342],order_in[338],order_in[334],order_in[330],order_in[326],order_in[322],order_in[318],order_in[314],order_in[310],order_in[306],order_in[302],order_in[298],order_in[294],order_in[290],order_in[286],order_in[282],order_in[278],order_in[274],order_in[270],order_in[266],order_in[262],order_in[258],order_in[254],order_in[250],order_in[246],order_in[242],order_in[238],order_in[234],order_in[230],order_in[226],order_in[222],order_in[218],order_in[214],order_in[210],order_in[206],order_in[202],order_in[198],order_in[194],order_in[190],order_in[186],order_in[182],order_in[178],order_in[174],order_in[170],order_in[166],order_in[162],order_in[158],order_in[154],order_in[150],order_in[146],order_in[142],order_in[138],order_in[134],order_in[130],order_in[126],order_in[122],order_in[118],order_in[114],order_in[110],order_in[106],order_in[102],order_in[98],order_in[94],order_in[90],order_in[86],order_in[82],order_in[78],order_in[74],order_in[70],order_in[66],order_in[62],order_in[58],order_in[54],order_in[50],order_in[46],order_in[42],order_in[38],order_in[34],order_in[30],order_in[26],order_in[22],order_in[18],order_in[14],order_in[10],order_in[6],order_in[2],order_in[357],order_in[353],order_in[349],order_in[345],order_in[341],order_in[337],order_in[333],order_in[329],order_in[325],order_in[321],order_in[317],order_in[313],order_in[309],order_in[305],order_in[301],order_in[297],order_in[293],order_in[289],order_in[285],order_in[281],order_in[277],order_in[273],order_in[269],order_in[265],order_in[261],order_in[257],order_in[253],order_in[249],order_in[245],order_in[241],order_in[237],order_in[233],order_in[229],order_in[225],order_in[221],order_in[217],order_in[213],order_in[209],order_in[205],order_in[201],order_in[197],order_in[193],order_in[189],order_in[185],order_in[181],order_in[177],order_in[173],order_in[169],order_in[165],order_in[161],order_in[157],order_in[153],order_in[149],order_in[145],order_in[141],order_in[137],order_in[133],order_in[129],order_in[125],order_in[121],order_in[117],order_in[113],order_in[109],order_in[105],order_in[101],order_in[97],order_in[93],order_in[89],order_in[85],order_in[81],order_in[77],order_in[73],order_in[69],order_in[65],order_in[61],order_in[57],order_in[53],order_in[49],order_in[45],order_in[41],order_in[37],order_in[33],order_in[29],order_in[25],order_in[21],order_in[17],order_in[13],order_in[9],order_in[5],order_in[1],order_in[356],order_in[352],order_in[348],order_in[344],order_in[340],order_in[336],order_in[332],order_in[328],order_in[324],order_in[320],order_in[316],order_in[312],order_in[308],order_in[304],order_in[300],order_in[296],order_in[292],order_in[288],order_in[284],order_in[280],order_in[276],order_in[272],order_in[268],order_in[264],order_in[260],order_in[256],order_in[252],order_in[248],order_in[244],order_in[240],order_in[236],order_in[232],order_in[228],order_in[224],order_in[220],order_in[216],order_in[212],order_in[208],order_in[204],order_in[200],order_in[196],order_in[192],order_in[188],order_in[184],order_in[180],order_in[176],order_in[172],order_in[168],order_in[164],order_in[160],order_in[156],order_in[152],order_in[148],order_in[144],order_in[140],order_in[136],order_in[132],order_in[128],order_in[124],order_in[120],order_in[116],order_in[112],order_in[108],order_in[104],order_in[100],order_in[96],order_in[92],order_in[88],order_in[84],order_in[80],order_in[76],order_in[72],order_in[68],order_in[64],order_in[60],order_in[56],order_in[52],order_in[48],order_in[44],order_in[40],order_in[36],order_in[32],order_in[28],order_in[24],order_in[20],order_in[16],order_in[12],order_in[8],order_in[4],order_in[0],order_in[359],order_in[355],order_in[351],order_in[347],order_in[343],order_in[339],order_in[335],order_in[331],order_in[327],order_in[323],order_in[319],order_in[315],order_in[311],order_in[307],order_in[303],order_in[299],order_in[295],order_in[291],order_in[287],order_in[283],order_in[279],order_in[275],order_in[271],order_in[267],order_in[263],order_in[259],order_in[255],order_in[251],order_in[247],order_in[243],order_in[239],order_in[235],order_in[231],order_in[227],order_in[223],order_in[219],order_in[215],order_in[211],order_in[207],order_in[203],order_in[199],order_in[195],order_in[191],order_in[187],order_in[183]};
			default:order_out <= 360'h00;
			endcase
		end
		else begin
			order_out <= 360'h00;
		end
	end
	else begin
	end
end

endmodule
