`timescale 1ns / 1ps
module F_normal_t12_next_Rom4(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b110100000011101001110100011110010011101010110011100001000101110010111100010001011000110111110110011011000100101010000000111110000001010100100000000101110000101110101101001110110111101100101001;
			5'h16: rd_q <= 192'b110010101110110100000000100000100110010011011111010001110101001101110111011100010111100111000101010101111010111110011010011001111110111110010001001101011111110111010011001100010010111100110111;
			5'h15: rd_q <= 192'b101111011000000100001100110001110100010010010010010100100110110100110110111111101101110011111101110111011011101101110010101011000001010100001000111000001111011001001100111110010101010111101000;
			5'h14: rd_q <= 192'b100110101011100001000101010111110011000111001111100111111101111010111101101111110000111000111001110110101100000001111110110011010010101101010010100011000111001111001011100100111010100101011001;
			5'h13: rd_q <= 192'b000010000001001000011010110000001100101101101001100111010110000001010010000001100001000111110100001001101000011001000001001100000010101100010110101101001000101100100010010101011111011000000101;
			5'h12: rd_q <= 192'b010010111111100011110110101100001100000100101100101000111000100010001101101111000101101001011010110010010100011110101010111000001011011000111101100100010101100001011000010001001001111000011011;
			5'h11: rd_q <= 192'b001111001100110111000111011011010110101000110101100111110100101100101011001001110111000111011101110111101000011101100110110110100000001111000011110111100101010011100010100010001111111111111000;
			5'h10: rd_q <= 192'b111101010001100101100001101010110011000111000101111101010010101111000001000010001001010000001110000101000011111110100101001111010000011000010000000111010001100110110001101010111110011001000100;
			5'h0f: rd_q <= 192'b111111001001011101000011000010001010111000011001000101000111101110101100011110110011010001001001101011101001111111110101010101100001001101011001001111001010100111101110111001000100000000111001;
			5'h0e: rd_q <= 192'b101001011110000111000101100010101011111101101111001000001111101100001010110010110000010011100110000001101001000110101000111101100001101011000011000101101000001010101001111001001100111010111011;
			5'h0d: rd_q <= 192'b000001011100100101001110010001111110101110100011101001000111100001111100111001000010110110001101101001001000010110001100000110101001101101001101101011100101101101001000001001010100011010110100;
			5'h0c: rd_q <= 192'b110110010111100001001011001100100010010011011111001101101100001011001001101000001110011001111001100010001000010011101101110111001111110111110111101010001101011011100100011011111101101100001011;
			5'h0b: rd_q <= 192'b010100110111111100101111111011110100001011110100101000011110011000111011110010010010111011111011000100110011101001000010011110010110010011011100010011100011100110110100101000101110101000001010;
			5'h0a: rd_q <= 192'b100101111011001010110110011110111110110010001101011000001000101000111101111001110111000110111000100000011101000101100011000000010111010101001001110100111001011110011111011110010011010100110000;
			5'h09: rd_q <= 192'b101100011111011100001010111101101000010110000001110110100010100001100101110000110010001111011110100010111000010011111001010011111110110010001001101001110010111011111110001001010011101011101100;
			5'h08: rd_q <= 192'b000101010000001101001001000000110111001011110110101011001011100000110111110111100101100100000110110101001000011111110010001100001111101010110001001111001001000000000100110011001010110011010000;
			5'h07: rd_q <= 192'b111110110100101000001011001000110011000100100111001010000011010000111011000001010110011111100101011111101000011011101010100110010100111101100001110011000101100101101001010110101010010001010000;
			5'h06: rd_q <= 192'b000111000000111000000010000001111111111011000101000110110111000000100110000110010001000011100000100001100001100000011000100010111101111001011110001001101000100001100001010001110101011000101010;
			5'h05: rd_q <= 192'b010010011011110100010111001010010101000001111000110010110100000000011110101011100010011010110011010001111011110110001110100100110011000101011011111001010101011010011111100000001010110111100010;
			5'h04: rd_q <= 192'b000011011010110110110000000100001101110000010100111000010110110001001011010010111110011001010101111011101001100000100001011100100001100001011011110100001010111111001101100011010100011101111011;
			5'h03: rd_q <= 192'b100100010001111001100010011001111110100110110001110011000001100100110010001111010101011101001001100000011100001100001111000111000011101110000000000100011010110001000100100010010111100101110110;
			5'h02: rd_q <= 192'b000010100100100001000001011001101010010111010000001001110111110100010110111011111111000001000101110011001000011111111000011010111100011010010101010110101000101000111001010111011100110110001100;
			5'h01: rd_q <= 192'b101110000010110100000110000001001100000101001111100101100101010110011111011100011010010011111101000111111010001101000111011111000111010001110110100010011101010011110001100111111001101101110000;
			5'h00: rd_q <= 192'b110000100000110110110101011101011000110101111100111010011011111011110010111010011110001100010110010000111000000011110010111011101000110111001101100001010110010001011101111100111110111001111011;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
