`timescale 1ns / 1ps
module F_normal_t12_next_Rom2(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b110111100100000011010000011111110101010001001001100110100111000010110101010101001000011100110101110111011111100111001111110010001011011010101000101101001010100110110001001011000111110101101110;
			5'h16: rd_q <= 192'b101101010001110100000011100100100010110111111010100101100100111110011001100001110101011111111001001100100110110110100101101101110101110001101100001111110111000001001001000001010010110100010110;
			5'h15: rd_q <= 192'b101001111111100110110010010010110111001110001101000001110011011110111101100110001001101101101101001011000101011111100000100011001100011100011111000111110001110110110100110001000000111010001111;
			5'h14: rd_q <= 192'b001110110001110010010100001010101010011011111010001100011111100110010000100111111101000001111101001100011011101111010001000010000011111001110110101011010000101110101001011011111111110001001011;
			5'h13: rd_q <= 192'b001000000100100001101011000000110010110110100110011101011000000101001000000110000100011111010000100110100001100100000100110000001010110001011010110100100010110010001001010101111101100000010100;
			5'h12: rd_q <= 192'b111000001011011101011010000011101101101111110001010010111010001100010100110100000011000100011101000100110111011101001101100101101010100111100010001100010010001011100011111100101011000010001001;
			5'h11: rd_q <= 192'b111100110011011100011101101101011010100011010110011111010010110010101100100111011100011101110111011110100001110110011011011010000000111100001111011110010101001110001010001000111111111111100000;
			5'h10: rd_q <= 192'b010010101100110010000111001101110111100110010000010111111010110101000000011000001110000011010100001111000010110101011000110111001111101001101000100111001110000111000011011011100000100011011010;
			5'h0f: rd_q <= 192'b011011001111010000001101101110010000011011100011110110101110110011110101101011100110000111001010110101101010110000011001011100001010111101001100000110100010000010111110010100001001000100101110;
			5'h0e: rd_q <= 192'b110001100111101010010111011111001001110001111000110011010110111101001101010011111111101100000010010000001111110010001001111001001111100000110000110001101100111000100000101100100110001111000011;
			5'h0d: rd_q <= 192'b000101110010010100111001000111111010111010001110100100011110000111110011100100001011011000110110100100100001011000110000011010100110110100110110101110010110110100100000100101010001101011010000;
			5'h0c: rd_q <= 192'b111110110100100000101101010100110010110111111011010100000000100101100010110000010010100100001010010011101100000001111011010110110001010111110110010010111101110010010100011111101111110111100110;
			5'h0b: rd_q <= 192'b100000101010100000111111011100001101010010010001010000100001100111001101000001011110001110011010011110101000000011101111111100011110001001100101010011001010010101010000011010110110000011001101;
			5'h0a: rd_q <= 192'b000011110011011101011000101110011101001111110001110011001010101110010001111111100010111001111000010111011111111110100110001110010100011000011011110100101001101011111010110001011000110111101111;
			5'h09: rd_q <= 192'b100101100010000110101010100011000111011111000011001001100010001011110001011011110110011111100000011101001010100111001111000000110010000100011010000000000111111101111111101101011011001010011111;
			5'h08: rd_q <= 192'b010101000000110100100100000011011100101111011010101100101110000011011111011110010110010000011011010100100001111111001000110000111110101011000100111100100100000000010011001100101011001101000000;
			5'h07: rd_q <= 192'b011100111000000100101101000101110111101000011011001010111101001010101000010101110010111101111001100101101100100001100110010011011101111110101111110110011110001010100000101010110000000010001010;
			5'h06: rd_q <= 192'b011100000011100000001000000111111111101100010100011011011100000010011000011001000100001110000010000110000110000001100010001011110111100101111000100110100010000110000101000111010101100010101000;
			5'h05: rd_q <= 192'b111010011010000011011100011010001001111010100000111010001000000101011000100110011100001010111011001010001001111111011100010110001011010001111011111000010001100111111100111000100111111101101101;
			5'h04: rd_q <= 192'b001101101011011011000000010000110111000001010011100001011011000100101101001011111001100101010111101110100110000010000101110010000110000101101111010000101011111100110110001101010001110111101100;
			5'h03: rd_q <= 192'b000101011000010000001000110010011100011100000011011111101110011110101110100101101011010110111100010111011011011000010110010011000111110100111100110110100111010110010101000001001011110011110111;
			5'h02: rd_q <= 192'b001010010010000100000101100110101001011101000000100111011111010001011011101111111100000100010111001100100001111111100001101011110001101001010101011010100010100011100101011101110011011000110000;
			5'h01: rd_q <= 192'b101100010100100110011001010001010110010011111010000101111101010100011011101001010111101101101110001001000011011100110111110011010100001011100110101110111001011101000001010111110011010011101111;
			5'h00: rd_q <= 192'b100101101001111111010100010011011000101101110100001011011111100110001111111001010011110010110101011000101101000000000111100100101101010100011110111111010001011001110010000011100010100000100110;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
