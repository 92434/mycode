`timescale 1ns / 1ps
module F_normal_t12_next_Rom3(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b011011110010000001101000001111111010101000100100110011010011100001011010101010100100001110011010111011101111110011100111111001000101101101010100010110100101010011011000100101100011111010110111;
			5'h16: rd_q <= 192'b010110101000111010000001110010010001011011111101010010110010011111001100110000111010101111111100100110010011011011010010110110111010111000110110000111111011100000100100100000101001011010001011;
			5'h15: rd_q <= 192'b101101000101011010011001010000110101011001100111011000010101101101001111110111001110000110001101100011010001111100000011010011000101101100000101101101011010111100011011000100100110001100110101;
			5'h14: rd_q <= 192'b111110100010010000001010011100111011110011011100111110100011110001011001010111110100010000000101100000111110100100011011100011100010011110110001011011001010010000010101110001111001101001010111;
			5'h13: rd_q <= 192'b000100000010010000110101100000011001011011010011001110101100000010100100000011000010001111101000010011010000110010000010011000000101011000101101011010010001011001000100101010111110110000001010;
			5'h12: rd_q <= 192'b100101111111000111101101011000011000001001011001010001110001000100011011011110001011010010110101100100101000111101010101110000010110110001111011001000101011000010110000100010010011110000110110;
			5'h11: rd_q <= 192'b011110011001101110001110110110101101010001101011001111101001011001010110010011101110001110111011101111010000111011001101101101000000011110000111101111001010100111000101000100011111111111110000;
			5'h10: rd_q <= 192'b001001010110011001000011100110111011110011001000001011111101011010100000001100000111000001101010000111100001011010101100011011100111110100110100010011100111000011100001101101110000010001101101;
			5'h0f: rd_q <= 192'b001101100111101000000110110111001000001101110001111011010111011001111010110101110011000011100101011010110101011000001100101110000101011110100110000011010001000001011111001010000100100010010111;
			5'h0e: rd_q <= 192'b100001001001011100001011110110001010000110011101100001000111011100110111101101110101000110111010001110110100101010110111111110000100010010010010010110010100011011010001001010010101010110010011;
			5'h0d: rd_q <= 192'b000010111001001010011100100011111101011101000111010010001111000011111001110010000101101100011011010010010000101100011000001101010011011010011011010111001011011010010000010010101000110101101000;
			5'h0c: rd_q <= 192'b011111011010010000010110101010011001011011111101101010000000010010110001011000001001010010000101001001110110000000111101101011011000101011111011001001011110111001001010001111110111111011110011;
			5'h0b: rd_q <= 192'b101001101111111001011111110111101000010111101001010000111100110001110111100100100101110111110110001001100111010010000100111100101100100110111000100111000111001101101001010001011101010000010100;
			5'h0a: rd_q <= 192'b111000000011000111101100001110100000011001011001000001001001010101011001111011111011101100000111001101011100101100100000000101101001101110000111110100110110110010111100000100101010001010000101;
			5'h09: rd_q <= 192'b101011001011101010010101001000001101010001000000011100011101000111101001101001110001111111001011001000010110000000010100100010111010100000000111001110100001111001111110101010101011110100111101;
			5'h08: rd_q <= 192'b001010100000011010010010000001101110010111101101010110010111000001101111101111001011001000001101101010010000111111100100011000011111010101100010011110010010000000001001100110010101100110100000;
			5'h07: rd_q <= 192'b001110011100000010010110100010111011110100001101100101011110100101010100001010111001011110111100110010110110010000110011001001101110111111010111111011001111000101010000010101011000000001000101;
			5'h06: rd_q <= 192'b001110000001110000000100000011111111110110001010001101101110000001001100001100100010000111000001000011000011000000110001000101111011110010111100010011010001000011000010100011101010110001010100;
			5'h05: rd_q <= 192'b100100110111101000101110010100101010000011110001100101101000000000111101010111000100110101100110100011110111101100011101001001100110001010110111110010101010110100111111000000010101101111000100;
			5'h04: rd_q <= 192'b000110110101101101100000001000011011100000101001110000101101100010010110100101111100110010101011110111010011000001000010111001000011000010110111101000010101111110011011000110101000111011110110;
			5'h03: rd_q <= 192'b111011010110100001000100000000100000110000100000010111011011001101000110010110111111011011100101001101011110111111111000001011000000011000010100010101110001101100001011111100100011101000001001;
			5'h02: rd_q <= 192'b000101001001000010000010110011010100101110100000010011101111101000101101110111111110000010001011100110010000111111110000110101111000110100101010101101010001010001110010101110111001101100011000;
			5'h01: rd_q <= 192'b101111110000111010001100110001000101110111011100111010010010101000011100110000100001000110001100000010010010111101101000111011001001100111111001011001111110101001100001110111111111111000000101;
			5'h00: rd_q <= 192'b010010110100111111101010001001101100010110111010000101101111110011000111111100101001111001011010101100010110100000000011110010010110101010001111011111101000101100111001000001110001010000010011;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
