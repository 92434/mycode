`timescale 1ns / 1ps
module F_normal_t12_next_Rom7(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[191:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 192'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h17: rd_q <= 192'b110001000100011110011110111100000111001100011111111010101111101100100010110111000011011010001011000100000111000010011111110101111011010000001100101101100100100011000100100010110001001000001011;
			5'h16: rd_q <= 192'b010100110110001000010000001110101000000010100011011000010011101000000010001000100101001000101011111000011010001010110110000010110110111110010101101101010010011100101010100000100000111011000011;
			5'h15: rd_q <= 192'b000101111011000000100001100110001110100010010010010010100100110110100110110111111101101110011111101110111011011101101110010101011000001010100001000111000001111011001001100111110010101010111101;
			5'h14: rd_q <= 192'b110011010001011111011000110101001011001001110000011010011000101101100010111000110110011011110010111001101010000111000000000100010001001111000010111001010010011111001000010111100000100001000101;
			5'h13: rd_q <= 192'b001110001110100011010011010000011010001010000101010010110001110000101110000001001110100100110000010000100001110111110100111001001000101101000000010110000001100100010100000101101010011111011100;
			5'h12: rd_q <= 192'b101001001110101011101110100110100011101110111100111111110110000111101100011010110101101001100011000010010100101101000011000100011011110000101010000110111001001001011010100111001101110010010100;
			5'h11: rd_q <= 192'b000001111001100110111000111011011010110101000110101100111110100101100101011001001110111000111011101110111101000011101100110110110100000001111000011110111100101010011100010100010001111111111111;
			5'h10: rd_q <= 192'b111110010000100101101100010100111000100110011001010111000110010111101001001100011011111010111010110110011011001100000111101011011001100001001000001110011000001011110111010001010001100010111010;
			5'h0f: rd_q <= 192'b110000011101001000111000000111100100000110001010101110001111111111000000110110111110000110111100111010000010101000110001011000100111010011000011100100110011110010001100111100001111010101101001;
			5'h0e: rd_q <= 192'b101110010010100111001000111111010111010001110100100011110000111110011100100001011011000110110100100100001011000110000011010100110110100110110101110010110110100100000100101010001101011010000000;
			5'h0d: rd_q <= 192'b111001110001001101101001101011100001001011010101100101100100111110011110100011000010100110001010101011111010010001000010100010010110101111100011100011111110101010101000011101001100110010100100;
			5'h0c: rd_q <= 192'b101101101011101011111001001010100110011100000010100011011100100010100100111010001100110111100111011000010111001100101011111101100011010101010011010111001010001110001101000110011011010000110110;
			5'h0b: rd_q <= 192'b011110011011101011000101110011101001111110001110011001010101110010001111111100010111001111000010111011111111110100110001110010100011000011011110100101001101011111010110001011000110111101111000;
			5'h0a: rd_q <= 192'b000100101111011001010110110011110111110110010001101011000001000101000111101111001110111000110111000100000011101000101100011000000010111010101001001110100111001011110011111011110010011010100110;
			5'h09: rd_q <= 192'b111100011001010010100001001110000011111100010001110110011000010110011101101010001100100001000000110010100100010001101100001000111100010100011011000011101100010000011110101101001100001100101111;
			5'h08: rd_q <= 192'b000000101010000001101001001000000110111001011110110101011001011100000110111110111100101100100000110110101001000011111110010001100001111101010110001001111001001000000000100110011001010110011010;
			5'h07: rd_q <= 192'b000111110110100101000001011001000110011000100100111001010000011010000111011000001010110011111100101011111101000011011101010100110010100111101100001110011000101100101101001010110101010010001010;
			5'h06: rd_q <= 192'b011100000101010011100000011100111000100000001000010100100000111001001100010010110111010000000001100111010101100101111010100101000110011110001110110110011100000111101100100100001101100011111100;
			5'h05: rd_q <= 192'b011110101110001010000010110101100101110111011111111010000000100001001011010111011001001011001011111001010110110111001000010101110111101001101110011000011011101000110011010010000010011110000101;
			5'h04: rd_q <= 192'b101011000010000001000110010011100011100000011011111101110011110101110100101101011010110111100010111011011011000010110010011000111110100111100110110100111010110010101000001001011110011110111000;
			5'h03: rd_q <= 192'b100001100101110010101100000110010110010101000111001010100010001111111111110111110101000011001111101001101001011011101011011011001010001110111111001001010000010010101001010110010111100101100101;
			5'h02: rd_q <= 192'b111001101110001101001000010010100011101100011011111001100010111100110011110011010101001000110011101000101010010000001100000001110100000001011000100100010111000010000110010110111101110111000011;
			5'h01: rd_q <= 192'b000101110000010110100000110000001001100000101001111100101100101010110011111011100011010010011111101000111111010001101000111011111000111010001110110100010011101010011110001100111111001101101110;
			5'h00: rd_q <= 192'b101101011101010001000110111000101001001000110110111101100010011100100011100000011110110101001010100110000001001110101000000100000111101101010100000110010001010111011010001010100011001010011000;
		default:rd_q <= 192'b0;
		endcase
	end
end

endmodule
