
`timescale 1ns / 1ps
module F_short_t12_next_Rom1(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[167:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 168'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h14: rd_q <= 168'b010100101101000001001100010001011111010111110011111110001010010101001011000001001110001011100010010110011010001100100110110010110000110010101011111011011010001100000001;
			5'h13: rd_q <= 168'b010000100101000011001010111011011000010111110010000001010001110001111101000100101000001100011101100000010110111011110010101010001001100001110101101011000100101011011110;
			5'h12: rd_q <= 168'b111100001000100100000010101000101000001101100001010110111010010110111111100110000101110010011100110000000011001100101110111101010101010111001011101000101111111001100001;
			5'h11: rd_q <= 168'b100111001110101001100001010011111000011001101001011000100000001000000101011010010100100111110100001110011100001110011010100110000011010110000101000011000011000100000000;
			5'h10: rd_q <= 168'b000000001001110011101010011000010100111110000110011010010110001000000010000001010110100101001001111101000011100111000011100110101001100000110101100001010000110000110001;
			5'h0f: rd_q <= 168'b100010001010111001100111101101100011100011011001011110110001100110010000000101011110110001111001011110101001111101011001110001111001100101100010000010010111111000110010;
			5'h0e: rd_q <= 168'b010011100010000001111010110110011010111110100110001111110010011010000011011011010111010011111101111011110100100000001101110011110011000111101000010101100001101111000111;
			5'h0d: rd_q <= 168'b011100100111000110000000110001100101000001100011100011011111101111011110000100010101011000100111010110000000001000001100110101110101000000001101011111100100101101101110;
			5'h0c: rd_q <= 168'b100111111011010101011010100111101101101011000010001100001111001111100100011111001111010001100010000110011111000000111110000101110110001111010111001110100011011000100001;
			5'h0b: rd_q <= 168'b110011100101010100010001010100100100111111000011001110011100110000011000001101100100111110111110100111101011100101111111010000111101101100011000111111010000101011001001;
			5'h0a: rd_q <= 168'b001100110010111000101100010111110010001111111100010011100011111001010011101001111011111001111111111000111110111100111001100001101111101111001001011110011001110010010110;
			5'h09: rd_q <= 168'b001001001011101010000111001000000110101110010100110111110100011101001100010110010010001110101010001011110101000100110011110111111000100110010100101000111010101101010100;
			5'h08: rd_q <= 168'b010101111101100111110010000001101000101011000111010100111111000001011000111110001111010111101111110101100001011001000101100101000110001111101000110001111101101010011010;
			5'h07: rd_q <= 168'b111000010000010110011100010011110100101001001101101011110101000001010101110011001100000001111100100000011001011010101101100111000001101011010000011110100010011100000001;
			5'h06: rd_q <= 168'b010000101110001100011111001111011000111101001101101110110100101110001000000011000100101100111111000111111011011011000111001000111100111101100011110101111101110101011010;
			5'h05: rd_q <= 168'b000101100110000001110010011011000110111101011100001011000101011100110011000100010001001111100100101110111011101001100110010000111011100010000000110001111101001000000101;
			5'h04: rd_q <= 168'b000000010101110100100001010000110111101110111000100100111100111011000010000111110000001010011000011011011101110100110110111111010110111110001010001011110111000101011110;
			5'h03: rd_q <= 168'b010101010110101010010111110000101100011001111000111000000111100111111011001011101001010011011001111101101001100111010000101001110001100101101011100001100011101101011000;
			5'h02: rd_q <= 168'b100100100111001111001110101001110001000000011010111101001100010110110001110100010011111011000101100110110011110111101010010010001001101010100100110000001100110100011001;
			5'h01: rd_q <= 168'b100000100110011010000001000110100100000000111000100110001001000010011110110001101010010001110010101111011100010000111001001101110010101011110101111001011000111110010011;
			5'h00: rd_q <= 168'b001001010100000010001110101111000011100100100000110101000111001101110111101110000101000100111011101010110110100110010100010001000001010001110111001100001000000111001011;
		default:rd_q <= 168'b0;
		endcase
	end
end

endmodule
