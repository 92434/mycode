
`timescale 1ns / 1ps
module F_short_t12_next_Rom2(
input	          							clk_1x,
input	          							rst_n,
//////////////////////////////////////////////////////////////
input										rd_en,
input				[4:0]				rdaddr,
output		reg			[167:0]				rd_q
);

always @(posedge clk_1x)begin
	if(~rst_n)begin
		rd_q <= 168'b0;
	end
	else if(rd_en == 1'b1)begin
		case(rdaddr)
			5'h14: rd_q <= 168'b100011001100100010111110101010010001000100011110000011010001100000110011100010111011010010110101100111111001011111011110111100111001111100000010001011011001011110000010;
			5'h13: rd_q <= 168'b001000010010100001100101011101101100001011111001000000101000111000111110100010010100000110001110110000001011011101111001010101000100110000111010110101100010010101101111;
			5'h12: rd_q <= 168'b110111011110010000011001110110101010101001010111010111001001100001001001110001011110101110001010110100110101111111011010111011001011001110110010000010100011100100110010;
			5'h11: rd_q <= 168'b010011100111010100110000101001111100001100110100101100010000000100000010101101001010010011111010000111001110000111001101010011000001101011000010100001100001100010000000;
			5'h10: rd_q <= 168'b101001011110111011101101101110110100110000100100110001011111101110010111000010110111000101100000010010010101101010101100010110110101010101001101000110011100000000011010;
			5'h0f: rd_q <= 168'b010001000101011100110011110110110001110001101100101111011000110011001000000010101111011000111100101111010100111110101100111000111100110010110001000001001011111100011001;
			5'h0e: rd_q <= 168'b100000101011000010100101111001110011110000110100111011101101100111010111101111110111111110111010010001001110001001001011011100011000000110100011111100000100101111100001;
			5'h0d: rd_q <= 168'b001110010011100011000000011000110010100000110001110001101111110111101111000010001010101100010011101011000000000100000110011010111010100000000110101111110010010110110111;
			5'h0c: rd_q <= 168'b111010100111101000110101110001001000011010000110111010010011001101100100001101111011111111110101101111111011111001010010100111011010100010111100010001100101110100010010;
			5'h0b: rd_q <= 168'b110000101000101000010000001000101100110000000110011011011010110010011010000100101110001000011011111111000001101011110010001101111111010011011011101001011100001101100110;
			5'h0a: rd_q <= 168'b000110011001011100010110001011111001000111111110001001110001111100101001110100111101111100111111111100011111011110011100110000110111110111100100101111001100111001001011;
			5'h09: rd_q <= 168'b000100100101110101000011100100000011010111001010011011111010001110100110001011001001000111010101000101111010100010011001111011111100010011001010010100011101010110101010;
			5'h08: rd_q <= 168'b001010111110110011111001000000110100010101100011101010011111100000101100011111000111101011110111111010110000101100100010110010100011000111110100011000111110110101001101;
			5'h07: rd_q <= 168'b110101010010001001010110101011000100111011000001001001101110001010111100111011111010010111111010111100111000110100011011010110000001010000111111111001100101010110000010;
			5'h06: rd_q <= 168'b001000010111000110001111100111101100011110100110110111011010010111000100000001100010010110011111100011111101101101100011100100011110011110110001111010111110111010101101;
			5'h05: rd_q <= 168'b101011101001000010100001101111011101110001001001111001110110000100001111100000010100110000110110111011101001101101111110101101111100010100010111101110001010111100000000;
			5'h04: rd_q <= 168'b000000001010111010010000101000011011110111011100010010011110011101100001000011111000000101001100001101101110111010011011011111101011011111000101000101111011100010101111;
			5'h03: rd_q <= 168'b001010101011010101001011111000010110001100111100011100000011110011111101100101110100101001101100111110110100110011101000010100111000110010110101110000110001110110101100;
			5'h02: rd_q <= 168'b111011001001100101111111110110000110001111101010100010110010100001001110111000010101101010100110011111101101100010111000101100100101010000000101101110110010000010001110;
			5'h01: rd_q <= 168'b111001001001001111011000000001101100101111111011101111010000001011011001011010101001011111111101111011011010010001010001000011011000110000101101001010011000000111001011;
			5'h00: rd_q <= 168'b101101110000000011011111110101011111011101110111100110110111001100101101110101011110110101011001011001101111001010000111101101000001001101101100010000110000011011100111;
		default:rd_q <= 168'b0;
		endcase
	end
end

endmodule
